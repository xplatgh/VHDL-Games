library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity bigbang is
port(
	clk,rst : in std_logic;
	rxd : in std_logic;
	hs,vs,r,g,b : out std_logic);
end bigbang;

architecture one of bigbang is

signal md : std_logic;
signal hs1,vs1,fclk,cclk,sclk : std_logic;
signal fs : std_logic_vector(2 downto 0);
signal cc : std_logic_vector(8 downto 0);
signal ll : std_logic_vector(8 downto 0);
signal grbx : std_logic_vector(3 downto 1);
signal grby : std_logic_vector(3 downto 1);
signal grbp : std_logic_vector(3 downto 1);
signal grb : std_logic_vector(3 downto 1);
signal grbc : std_logic_vector(3 downto 1);
signal mode : std_logic_vector(2 downto 0);

signal clk_cnt,clk_rsclk : std_logic_vector(24 downto 0);
signal PT0,PT1,PT2,PT3,PT4,PT5 : std_logic_vector(3 downto 0);
signal pt : std_logic;

signal freq,scal, sin,tri,squ,rl : std_logic;
type index_type is array(0 to 800) of integer range 0 to 200;
signal tri_ind,squ_ind,sin_ind,sin_id : index_type;
signal x : integer range 0 to 200;
signal sin_y,tri_y,squ_y : integer range 0 to 200;
signal wi : integer range 0 to 7;
signal f,sc,rlf : integer range 1 to 8;
signal cci : integer range 0 to 511;
signal rrll : integer range 0 to 200;
signal xt,xf : integer range 0 to 1800;

signal clk_rscnt:integer range 0 to 651;
signal sam_clk:std_logic;
signal done : std_logic;
type status_type is(start,data,over);
signal status:status_type;
signal sam_cnt:std_logic_vector(2 downto 0);
signal bit_cnt:std_logic_vector(3 downto 0);
signal rcv_shift_reg:std_logic_vector(7 downto 0);
signal rcv_data:std_logiC_vector(7 downto 0);
signal rrr,l,rot,rev,speed,pul : std_logic;
signal rrrr,uu,lll,dd : std_logic;

type status_stype is array(0 to 17,0 to 17) of std_logic;    --(250-2*2)*(400-4*2)/8=12054--------------64x64--------------
type index_stype is array(0 to 100) of integer range 0 to 127;       --max : 12054--------------4096-------
signal status1,status0 : status_stype;
signal index_x,index_y : index_stype;
signal alive : std_logic;
signal di,dir : std_logic_vector(1 downto 0);
signal i,j,k,m,n : integer range 0 to 127;
signal len : integer range 0 to 100;
signal food : std_logic;
signal food_x,food_y : integer range 1 to 16;
signal lcx : std_logic;
signal score1,score0 : std_logic_vector(3 downto 0);
signal ccc,llc : integer range 0 to 127;

type ttstatus_type is array(0 to 11,0 to 42) of std_logic;    --(250-2*2)*(400-4*2)/8=12054
type index_typex is array(0 to 3) of integer range 0 to 15;
type index_typey is array(0 to 3) of integer range 0 to 63;
type tstatuse_type is (start,usual,dead);
signal ttstatus1,ttstatus0 : ttstatus_type;
signal tindex_x : index_typex;
signal tindex_y : index_typey;
signal tstatus : tstatuse_type;
signal food0,food1 : integer range 0 to 6;
signal tra,tra_r,tra_l,tra_ro,tra_re,tra_d : std_logic;
signal ti,tj,tk,tm,tn,tsp : integer range 0 to 63;
signal tccc,tlll : integer range 0 to 511;

begin
grb(2)<=(grbp(2))and hs1 and vs1;
grb(3)<=(grbp(3))and hs1 and vs1;
grb(1)<=(grbp(1))and hs1 and vs1;

process(clk)
begin
if rising_edge(clk) then
if (md='1') then
end if;
end if;
end process;

------------------------------------rs232-------------------------------

P1:process(clk,rst)
begin
	if rst='0' then
		clk_rscnt<=0;
	elsif rising_edge(clk) then
		if clk_rscnt=651 then
			clk_rscnt<=0;
			sam_clk<='1';
		else
			clk_rscnt<=clk_rscnt+1;
			sam_clk<='0';
		end if;
	end if;
end process P1;

P2:process(clk,rst)
begin
	if rst='0' then
		status<=start;
		sam_cnt<="000";
		bit_cnt<="0000";
		rcv_shift_reg<="00111111";
		rcv_data<="00111111";
		done<='1';

		freq<='0';
		scal<='0'; 
		sin<='1';
		tri<='1';
		squ<='1';
		rl<='0';
		rrll<=0;

		rrr<='0';
		l<='0';
		rot<='0';
		rev<='0';
		speed<='0';
		pul<='0';

		rrrr<='0';
		uu<='0';
		lll<='0';
		dd<='0';

	elsif rising_edge(clk) then
		if sam_clk='1' then
			case status is
				when start=>
					if rxd='0' then
						if sam_cnt="011" then
							sam_cnt<="000";
							status<=data;
							bit_cnt<="0000";
						else
							sam_cnt<=sam_cnt+'1';
						end if;
					end if;
				when data=>
					if sam_cnt="111" then
						if bit_cnt="1000" then
							status<=over;
						else
							rcv_shift_reg<=rxd&rcv_shift_reg(7 downto 1);
							sam_cnt<="000";
							bit_cnt<=bit_cnt+'1';
						end if;
					else
						sam_cnt<=sam_cnt+'1';
					end if;
				when over=>
					rcv_data<=rcv_shift_reg;
					if done='1' then
					if rcv_data="00001010" then
						if mode="111" then               
							mode<="000";
						else
							mode<=mode+1;
						end if;		
					end if;	
	
					if mode="101" then
						if rcv_data="01110001" then
							if f=8 then
							f<=1;
							else
							f<=f+1;
							end if;
						elsif rcv_data="01110111" then
							if sc=8 then
								sc<=1;
							elsif (sc=1 or sc=2 or sc=4) then
								sc<=sc*2;
							else
								sc<=1;
							end if;
							rlf<=sc;
						elsif rcv_data="01100101" then
							sin<=not sin;
						elsif rcv_data="01110010" then
							tri<=not tri;
						elsif rcv_data="01110100" then
							squ<=not squ;
						elsif rcv_data="01111001" then
							if rrll=200 then
								rrll<=0;
								if rlf=1 then
									rlf<=sc;
								else
									rlf<=rlf-1;
								end if;
							else 
								rrll<=rrll+1;
							end if;
						end if;			
					elsif mode="111" then
						if rcv_data="01100001" then
							rrr<=not rrr;
						elsif rcv_data="01110011" then
							l<=not l;
						elsif rcv_data="01100100" then
							rot<=not rot;
						elsif rcv_data="01100110" then
							rev<=not rev;
						elsif rcv_data="01100111" then
							speed<=not speed;
						elsif rcv_data="01101000" then
							pul<=not pul;
						end if;
					elsif mode="110" then
						if rcv_data="01111010" then
							rrrr<=not rrrr;
						elsif rcv_data="01111000" then
							uu<=not uu;
						elsif rcv_data="01100011" then
							lll<=not lll;
						elsif rcv_data="01110110" then
							dd<=not dd;
						end if;
					end if;
					end if;
					done<=not done;
					status<=start;
			end case;
		end if;
	end if;
end process P2;



    PROCESS( CLK )
    BEGIN
        IF CLK'EVENT AND CLK = '1' THEN -- 50MHz 5��Ƶ
            IF FS = 4 THEN FS <= "000";
            ELSE
                FS <= (FS + 1);
            END IF;
        END IF;
    END PROCESS;
    FCLK <= FS(2);
    PROCESS( FCLK )--��315��Ƶ��12000000/(13*30)=30769,�ӽ�����Ƶ31469
    BEGIN
        IF FCLK'EVENT AND FCLK = '1' THEN
            IF CC = 314 THEN  CC <= "000000000";
            ELSE
                CC <= CC + 1;
            END IF;
        END IF;
    END PROCESS;
    CCLK <= CC(8);
    
    PROCESS( CCLK )
    BEGIN
        IF CCLK'EVENT AND CCLK = '0' THEN
            IF LL = 481 THEN  LL <= "000000000";
            ELSE
                LL <= LL + 1;
            END IF;
        END IF;
    END PROCESS;
    
    
    PROCESS( CC,LL )
    BEGIN
        IF CC > 251 THEN  HS1 <= '0';  --��ͬ��
        ELSE
            HS1 <= '1';
        END IF;
        IF LL > 479 THEN  VS1 <= '0'; --��ͬ��
        ELSE
            VS1 <= '1';
        END IF;
    END PROCESS;
    
process(clk)
begin
	if rising_edge(clk) then
		IF clk_cnt=25000000 THEN clk_cnt<=(others=>'0');
        ELSE
            clk_cnt<=clk_cnt+1;
        END IF;
    END IF;
END PROCESS;

sclk<=clk_cnt(24);
----------------------------------------clk------------------------------
process(sclk,rst)
begin
if rst='0' then

PT0<="0000";PT1<="0000";PT2<="0000";PT3<="0000";PT4<="0000";PT5<="0000";pt<='0';

elsif rising_edge(sclk) then
pt<=not pt;
if pt='1' then
	if PT4="0101" and PT5="1001" then
		if PT2="0101" and PT3="1001" then
			if PT0="0010" and PT1="0011" then
				PT0<="0000";PT1<="0000";PT2<="0000";PT3<="0000";PT4<="0000";PT5<="0000";
			elsif PT1="1001" then
				PT0<=PT0+1;PT1<="0000";
			else
				PT1<=PT1+1;
			end if;
		elsif PT3="1001" then
			PT2<=PT2+1;PT3<="0000";
		else
			PT3<=PT3+1;
		end if;
	elsif PT5="1001" then
		PT4<=PT4+1;PT5<="0000";
	else
		PT5<=PT5+1;
	end if;
end if;
end if;
end process;

 ------------------------------------------wave--------------------------------- 
process(clk)
begin
if rising_edge(clk) then
	if x=200 then
		x<=0;
	else
		x<=x+1;
	end if;
end if;
end process;  

process(clk)
begin
if mode="101" then

	sin_ind(0)<=100;
	sin_ind(1)<=103;
	sin_ind(2)<=106;
	sin_ind(3)<=109;
	sin_ind(4)<=113;
	sin_ind(5)<=116;
	sin_ind(6)<=119;
	sin_ind(7)<=122;
	sin_ind(8)<=125;
	sin_ind(9)<=128;
	sin_ind(10)<=131;
	sin_ind(11)<=134;
	sin_ind(12)<=137;
	sin_ind(13)<=140;
	sin_ind(14)<=143;
	sin_ind(15)<=145;
	sin_ind(16)<=148;
	sin_ind(17)<=151;
	sin_ind(18)<=154;
	sin_ind(19)<=156;
	sin_ind(20)<=159;
	sin_ind(21)<=161;
	sin_ind(22)<=164;
	sin_ind(23)<=166;
	sin_ind(24)<=168;
	sin_ind(25)<=171;
	sin_ind(26)<=173;
	sin_ind(27)<=175;
	sin_ind(28)<=177;
	sin_ind(29)<=179;
	sin_ind(30)<=181;
	sin_ind(31)<=183;
	sin_ind(32)<=184;
	sin_ind(33)<=186;
	sin_ind(34)<=188;
	sin_ind(35)<=189;
	sin_ind(36)<=190;
	sin_ind(37)<=192;
	sin_ind(38)<=193;
	sin_ind(39)<=194;
	sin_ind(40)<=195;
	sin_ind(41)<=196;
	sin_ind(42)<=197;
	sin_ind(43)<=198;
	sin_ind(44)<=198;
	sin_ind(45)<=199;
	sin_ind(46)<=199;
	sin_ind(47)<=200;
	sin_ind(48)<=200;
	sin_ind(49)<=200;
	sin_ind(50)<=200;
	sin_ind(51)<=200;
	sin_ind(52)<=200;
	sin_ind(53)<=200;
	sin_ind(54)<=199;
	sin_ind(55)<=199;
	sin_ind(56)<=198;
	sin_ind(57)<=198;
	sin_ind(58)<=197;
	sin_ind(59)<=196;
	sin_ind(60)<=195;
	sin_ind(61)<=194;
	sin_ind(62)<=193;
	sin_ind(63)<=192;
	sin_ind(64)<=191;
	sin_ind(65)<=189;
	sin_ind(66)<=188;
	sin_ind(67)<=186;
	sin_ind(68)<=184;
	sin_ind(69)<=183;
	sin_ind(70)<=181;
	sin_ind(71)<=179;
	sin_ind(72)<=177;
	sin_ind(73)<=175;
	sin_ind(74)<=173;
	sin_ind(75)<=171;
	sin_ind(76)<=169;
	sin_ind(77)<=166;
	sin_ind(78)<=164;
	sin_ind(79)<=161;
	sin_ind(80)<=159;
	sin_ind(81)<=156;
	sin_ind(82)<=154;
	sin_ind(83)<=151;
	sin_ind(84)<=148;
	sin_ind(85)<=146;
	sin_ind(86)<=143;
	sin_ind(87)<=140;
	sin_ind(88)<=137;
	sin_ind(89)<=134;
	sin_ind(90)<=131;
	sin_ind(91)<=128;
	sin_ind(92)<=125;
	sin_ind(93)<=122;
	sin_ind(94)<=119;
	sin_ind(95)<=116;
	sin_ind(96)<=113;
	sin_ind(97)<=110;
	sin_ind(98)<=106;
	sin_ind(99)<=103;
	sin_ind(100)<=100;
	sin_ind(101)<=97;
	sin_ind(102)<=94;
	sin_ind(103)<=91;
	sin_ind(104)<=88;
	sin_ind(105)<=85;
	sin_ind(106)<=81;
	sin_ind(107)<=78;
	sin_ind(108)<=75;
	sin_ind(109)<=72;
	sin_ind(110)<=69;
	sin_ind(111)<=66;
	sin_ind(112)<=63;
	sin_ind(113)<=60;
	sin_ind(114)<=58;
	sin_ind(115)<=55;
	sin_ind(116)<=52;
	sin_ind(117)<=49;
	sin_ind(118)<=47;
	sin_ind(119)<=44;
	sin_ind(120)<=41;
	sin_ind(121)<=39;
	sin_ind(122)<=36;
	sin_ind(123)<=34;
	sin_ind(124)<=32;
	sin_ind(125)<=29;
	sin_ind(126)<=27;
	sin_ind(127)<=25;
	sin_ind(128)<=23;
	sin_ind(129)<=21;
	sin_ind(130)<=19;
	sin_ind(131)<=17;
	sin_ind(132)<=16;
	sin_ind(133)<=14;
	sin_ind(134)<=12;
	sin_ind(135)<=11;
	sin_ind(136)<=10;
	sin_ind(137)<=8;
	sin_ind(138)<=7;
	sin_ind(139)<=6;
	sin_ind(140)<=5;
	sin_ind(141)<=4;
	sin_ind(142)<=3;
	sin_ind(143)<=2;
	sin_ind(144)<=2;
	sin_ind(145)<=1;
	sin_ind(146)<=1;
	sin_ind(147)<=0;
	sin_ind(148)<=0;
	sin_ind(149)<=0;
	sin_ind(150)<=0;
	sin_ind(151)<=0;
	sin_ind(152)<=0;
	sin_ind(153)<=0;
	sin_ind(154)<=1;
	sin_ind(155)<=1;
	sin_ind(156)<=2;
	sin_ind(157)<=2;
	sin_ind(158)<=3;
	sin_ind(159)<=4;
	sin_ind(160)<=5;
	sin_ind(161)<=6;
	sin_ind(162)<=7;
	sin_ind(163)<=8;
	sin_ind(164)<=9;
	sin_ind(165)<=11;
	sin_ind(166)<=12;
	sin_ind(167)<=14;
	sin_ind(168)<=15;
	sin_ind(169)<=17;
	sin_ind(170)<=19;
	sin_ind(171)<=21;
	sin_ind(172)<=23;
	sin_ind(173)<=25;
	sin_ind(174)<=27;
	sin_ind(175)<=29;
	sin_ind(176)<=31;
	sin_ind(177)<=34;
	sin_ind(178)<=36;
	sin_ind(179)<=38;
	sin_ind(180)<=41;
	sin_ind(181)<=44;
	sin_ind(182)<=46;
	sin_ind(183)<=49;
	sin_ind(184)<=52;
	sin_ind(185)<=54;
	sin_ind(186)<=57;
	sin_ind(187)<=60;
	sin_ind(188)<=63;
	sin_ind(189)<=66;
	sin_ind(190)<=69;
	sin_ind(191)<=72;
	sin_ind(192)<=75;
	sin_ind(193)<=78;
	sin_ind(194)<=81;
	sin_ind(195)<=84;
	sin_ind(196)<=87;
	sin_ind(197)<=90;
	sin_ind(198)<=93;
	sin_ind(199)<=97;
	sin_ind(200)<=100;

if rising_edge(clk) then

if x>=rrll and rlf=sc then
	xf<=(x-rrll)*f/sc;
else
	xf<=(x+200*rlf-rrll)*f/sc;
end if;

for wi in  0 to 7 loop
	if xf>=200*wi and xf<200*(wi+1) then
		xt<=xf-200*wi;
	end if;
end loop;
	if xt<50 then
		tri_y<=100-xt*2;
	elsif xt<150 then
		tri_y<=(xt-50)*2;
	else
		tri_y<=200-(xt-150)*2;
	end if;
	if xt<100 then
		squ_y<=200;
	else
		squ_y<=0;
	end if;
		
	sin_id(x)<=sin_ind(xt);
	
tri_ind(x)<=tri_y;
squ_ind(x)<=squ_y;
end if;
end if;
end process;
		
---------------------snake------------------------

				
process(cc,ll)
begin 
	grbp<="000";


--------------------------------mode="000"--------------------vertical--------------------
if mode="000" or mode="010" then
 
if cc<31 then grby<="000";
end if;
if cc>=31 and cc<62 then grby<="001";
end if;
if cc>=62 and cc<93 then grby<="010";
end if;
if cc>=93 and cc<124 then grby<="011";
end if;
if cc>=124 and cc<155 then grby<="100";
end if;
if cc>=155 and cc<186 then grby<="101";
end if;
if cc>=186 and cc<217 then grby<="110";  
end if;
if cc>=217 and cc<251 then grby<="111";
end if; 
    
end if;

if mode="000" then
    grbp<=grby;
end if;


--------------------------------mode="001"------------------horizontal------------------
if mode="001" or mode="010" then

if ll<53 then grbx<="000";
end if;
if ll>=53 and ll<106 then grbx<="001";
end if;
if ll>=106 and ll<159 then grbx<="010";
end if;
if ll>=159 and ll<212 then grbx<="011";
end if;
if ll>=212 and ll<265 then grbx<="100";
end if;
if ll>=265 and ll<318 then grbx<="101";
end if;
if ll>=318 and ll<371 then grbx<="110";
end if;
if ll>=371 and ll<426 then grbx<="111";
end if;   
    
end if;

if mode="001" then
    grbp<=grbx;
end if;

--------------------------------mode="010"-------------------cross-------------------
if mode="010" then
    
grbc<=grbx xor grby;
if grbc(1)='0' then
    grbp<="111";
else
    grbp<="000";
end if;

end if;

-------------------------------mode="011"--------------------pic----------------------
if mode="011" then
	if (cc=13 and ll=0) then grbp<="010";
	end if;
	if (cc=27 and ll=0) then grbp<="010";
	end if;
	if (ll=0 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=0 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=0) then grbp<="010";
	end if;
	if (cc=183 and ll=0) then grbp<="010";
	end if;
	if (ll=0 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=0 and cc>=207 and cc<248) then grbp<="010";
	end if;
	if (cc=13 and ll=1) then grbp<="010";
	end if;
	if (cc=27 and ll=1) then grbp<="010";
	end if;
	if (ll=1 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=1 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=1) then grbp<="010";
	end if;
	if (cc=183 and ll=1) then grbp<="010";
	end if;
	if (ll=1 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=1 and cc>=207 and cc<248) then grbp<="010";
	end if;
	if (cc=13 and ll=2) then grbp<="010";
	end if;
	if (cc=27 and ll=2) then grbp<="010";
	end if;
	if (ll=2 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=2 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=2) then grbp<="010";
	end if;
	if (cc=183 and ll=2) then grbp<="010";
	end if;
	if (ll=2 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=2 and cc>=207 and cc<248) then grbp<="010";
	end if;
	if (cc=13 and ll=3) then grbp<="010";
	end if;
	if (cc=27 and ll=3) then grbp<="010";
	end if;
	if (ll=3 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=3 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=3) then grbp<="010";
	end if;
	if (cc=183 and ll=3) then grbp<="010";
	end if;
	if (ll=3 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=3 and cc>=207 and cc<248) then grbp<="010";
	end if;
	if (cc=6 and ll=4) then grbp<="010";
	end if;
	if (cc=10 and ll=4) then grbp<="010";
	end if;
	if (ll=4 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (cc=16 and ll=4) then grbp<="010";
	end if;
	if (cc=27 and ll=4) then grbp<="010";
	end if;
	if (ll=4 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=4 and cc>=168 and cc<170) then grbp<="010";
	end if;
	if (ll=4 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (cc=180 and ll=4) then grbp<="010";
	end if;
	if (ll=4 and cc>=180 and cc<186) then grbp<="010";
	end if;
	if (cc=196 and ll=4) then grbp<="010";
	end if;
	if (cc=207 and ll=4) then grbp<="010";
	end if;
	if (ll=4 and cc>=207 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=5) then grbp<="010";
	end if;
	if (cc=9 and ll=5) then grbp<="010";
	end if;
	if (ll=5 and cc>=9 and cc<12) then grbp<="010";
	end if;
	if (cc=27 and ll=5) then grbp<="010";
	end if;
	if (ll=5 and cc>=27 and cc<164) then grbp<="010";
	end if;
	if (ll=5 and cc>=169 and cc<173) then grbp<="010";
	end if;
	if (cc=179 and ll=5) then grbp<="010";
	end if;
	if (ll=5 and cc>=179 and cc<183) then grbp<="010";
	end if;
	if (ll=5 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (cc=208 and ll=5) then grbp<="010";
	end if;
	if (ll=5 and cc>=208 and cc<250) then grbp<="010";
	end if;
	if (ll=6 and cc>=7 and cc<9) then grbp<="010";
	end if;
	if (cc=13 and ll=6) then grbp<="010";
	end if;
	if (ll=6 and cc>=13 and cc<16) then grbp<="010";
	end if;
	if (ll=6 and cc>=27 and cc<163) then grbp<="010";
	end if;
	if (ll=6 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=6 and cc>=176 and cc<178) then grbp<="010";
	end if;
	if (cc=185 and ll=6) then grbp<="010";
	end if;
	if (cc=187 and ll=6) then grbp<="010";
	end if;
	if (cc=197 and ll=6) then grbp<="010";
	end if;
	if (cc=208 and ll=6) then grbp<="010";
	end if;
	if (ll=6 and cc>=208 and cc<248) then grbp<="010";
	end if;
	if (cc=11 and ll=7) then grbp<="010";
	end if;
	if (cc=14 and ll=7) then grbp<="010";
	end if;
	if (cc=16 and ll=7) then grbp<="010";
	end if;
	if (cc=27 and ll=7) then grbp<="010";
	end if;
	if (ll=7 and cc>=27 and cc<165) then grbp<="010";
	end if;
	if (cc=183 and ll=7) then grbp<="010";
	end if;
	if (cc=186 and ll=7) then grbp<="010";
	end if;
	if (cc=197 and ll=7) then grbp<="010";
	end if;
	if (cc=208 and ll=7) then grbp<="010";
	end if;
	if (ll=7 and cc>=208 and cc<248) then grbp<="010";
	end if;
	if (cc=7 and ll=8) then grbp<="010";
	end if;
	if (cc=11 and ll=8) then grbp<="010";
	end if;
	if (ll=8 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (cc=27 and ll=8) then grbp<="010";
	end if;
	if (ll=8 and cc>=27 and cc<165) then grbp<="010";
	end if;
	if (cc=172 and ll=8) then grbp<="010";
	end if;
	if (cc=187 and ll=8) then grbp<="010";
	end if;
	if (ll=8 and cc>=187 and cc<189) then grbp<="010";
	end if;
	if (cc=194 and ll=8) then grbp<="010";
	end if;
	if (cc=197 and ll=8) then grbp<="010";
	end if;
	if (cc=209 and ll=8) then grbp<="010";
	end if;
	if (ll=8 and cc>=209 and cc<247) then grbp<="010";
	end if;
	if (cc=9 and ll=9) then grbp<="010";
	end if;
	if (cc=11 and ll=9) then grbp<="010";
	end if;
	if (ll=9 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=9 and cc>=14 and cc<16) then grbp<="010";
	end if;
	if (ll=9 and cc>=27 and cc<166) then grbp<="010";
	end if;
	if (ll=9 and cc>=187 and cc<189) then grbp<="010";
	end if;
	if (ll=9 and cc>=190 and cc<192) then grbp<="010";
	end if;
	if (cc=197 and ll=9) then grbp<="010";
	end if;
	if (ll=9 and cc>=197 and cc<199) then grbp<="010";
	end if;
	if (ll=9 and cc>=209 and cc<246) then grbp<="010";
	end if;
	if (cc=13 and ll=10) then grbp<="010";
	end if;
	if (cc=27 and ll=10) then grbp<="010";
	end if;
	if (ll=10 and cc>=27 and cc<166) then grbp<="010";
	end if;
	if (cc=191 and ll=10) then grbp<="010";
	end if;
	if (ll=10 and cc>=191 and cc<193) then grbp<="010";
	end if;
	if (ll=10 and cc>=197 and cc<199) then grbp<="010";
	end if;
	if (ll=10 and cc>=209 and cc<246) then grbp<="010";
	end if;
	if (cc=27 and ll=11) then grbp<="010";
	end if;
	if (ll=11 and cc>=27 and cc<166) then grbp<="010";
	end if;
	if (cc=189 and ll=11) then grbp<="010";
	end if;
	if (cc=191 and ll=11) then grbp<="010";
	end if;
	if (ll=11 and cc>=191 and cc<193) then grbp<="010";
	end if;
	if (ll=11 and cc>=196 and cc<200) then grbp<="010";
	end if;
	if (ll=11 and cc>=210 and cc<245) then grbp<="010";
	end if;
	if (cc=27 and ll=12) then grbp<="010";
	end if;
	if (ll=12 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=12) then grbp<="010";
	end if;
	if (ll=12 and cc>=190 and cc<194) then grbp<="010";
	end if;
	if (cc=198 and ll=12) then grbp<="010";
	end if;
	if (ll=12 and cc>=198 and cc<200) then grbp<="010";
	end if;
	if (ll=12 and cc>=210 and cc<245) then grbp<="010";
	end if;
	if (cc=27 and ll=13) then grbp<="010";
	end if;
	if (ll=13 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (ll=13 and cc>=186 and cc<189) then grbp<="010";
	end if;
	if (cc=193 and ll=13) then grbp<="010";
	end if;
	if (cc=195 and ll=13) then grbp<="010";
	end if;
	if (ll=13 and cc>=195 and cc<200) then grbp<="010";
	end if;
	if (ll=13 and cc>=211 and cc<244) then grbp<="010";
	end if;
	if (cc=8 and ll=14) then grbp<="010";
	end if;
	if (cc=10 and ll=14) then grbp<="010";
	end if;
	if (cc=12 and ll=14) then grbp<="010";
	end if;
	if (ll=14 and cc>=12 and cc<14) then grbp<="010";
	end if;
	if (ll=14 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=188 and ll=14) then grbp<="010";
	end if;
	if (cc=191 and ll=14) then grbp<="010";
	end if;
	if (cc=193 and ll=14) then grbp<="010";
	end if;
	if (cc=195 and ll=14) then grbp<="010";
	end if;
	if (ll=14 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (ll=14 and cc>=211 and cc<243) then grbp<="010";
	end if;
	if (cc=26 and ll=15) then grbp<="010";
	end if;
	if (ll=15 and cc>=26 and cc<166) then grbp<="010";
	end if;
	if (cc=190 and ll=15) then grbp<="010";
	end if;
	if (cc=192 and ll=15) then grbp<="010";
	end if;
	if (cc=194 and ll=15) then grbp<="010";
	end if;
	if (ll=15 and cc>=194 and cc<196) then grbp<="010";
	end if;
	if (ll=15 and cc>=197 and cc<201) then grbp<="010";
	end if;
	if (ll=15 and cc>=211 and cc<243) then grbp<="010";
	end if;
	if (cc=12 and ll=16) then grbp<="010";
	end if;
	if (cc=27 and ll=16) then grbp<="010";
	end if;
	if (ll=16 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=16) then grbp<="010";
	end if;
	if (cc=192 and ll=16) then grbp<="010";
	end if;
	if (ll=16 and cc>=192 and cc<195) then grbp<="010";
	end if;
	if (ll=16 and cc>=196 and cc<201) then grbp<="010";
	end if;
	if (ll=16 and cc>=212 and cc<242) then grbp<="010";
	end if;
	if (cc=12 and ll=17) then grbp<="010";
	end if;
	if (cc=27 and ll=17) then grbp<="010";
	end if;
	if (ll=17 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=17) then grbp<="010";
	end if;
	if (ll=17 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (ll=17 and cc>=196 and cc<202) then grbp<="010";
	end if;
	if (ll=17 and cc>=212 and cc<241) then grbp<="010";
	end if;
	if (cc=26 and ll=18) then grbp<="010";
	end if;
	if (ll=18 and cc>=26 and cc<167) then grbp<="010";
	end if;
	if (cc=188 and ll=18) then grbp<="010";
	end if;
	if (cc=190 and ll=18) then grbp<="010";
	end if;
	if (ll=18 and cc>=190 and cc<202) then grbp<="010";
	end if;
	if (ll=18 and cc>=212 and cc<241) then grbp<="010";
	end if;
	if (cc=10 and ll=19) then grbp<="010";
	end if;
	if (cc=27 and ll=19) then grbp<="010";
	end if;
	if (ll=19 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=19) then grbp<="010";
	end if;
	if (cc=192 and ll=19) then grbp<="010";
	end if;
	if (cc=195 and ll=19) then grbp<="010";
	end if;
	if (ll=19 and cc>=195 and cc<202) then grbp<="010";
	end if;
	if (ll=19 and cc>=213 and cc<240) then grbp<="010";
	end if;
	if (ll=20 and cc>=1 and cc<3) then grbp<="010";
	end if;
	if (ll=20 and cc>=26 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=20) then grbp<="010";
	end if;
	if (ll=20 and cc>=190 and cc<196) then grbp<="010";
	end if;
	if (ll=20 and cc>=197 and cc<203) then grbp<="010";
	end if;
	if (ll=20 and cc>=213 and cc<240) then grbp<="010";
	end if;
	if (cc=26 and ll=21) then grbp<="010";
	end if;
	if (ll=21 and cc>=26 and cc<167) then grbp<="010";
	end if;
	if (cc=188 and ll=21) then grbp<="010";
	end if;
	if (ll=21 and cc>=188 and cc<193) then grbp<="010";
	end if;
	if (ll=21 and cc>=194 and cc<203) then grbp<="010";
	end if;
	if (ll=21 and cc>=213 and cc<239) then grbp<="010";
	end if;
	if (ll=22 and cc>=26 and cc<167) then grbp<="010";
	end if;
	if (cc=190 and ll=22) then grbp<="010";
	end if;
	if (ll=22 and cc>=190 and cc<192) then grbp<="010";
	end if;
	if (cc=197 and ll=22) then grbp<="010";
	end if;
	if (ll=22 and cc>=197 and cc<203) then grbp<="010";
	end if;
	if (ll=22 and cc>=214 and cc<238) then grbp<="010";
	end if;
	if (ll=23 and cc>=27 and cc<167) then grbp<="010";
	end if;
	if (cc=194 and ll=23) then grbp<="010";
	end if;
	if (ll=23 and cc>=194 and cc<198) then grbp<="010";
	end if;
	if (ll=23 and cc>=199 and cc<204) then grbp<="010";
	end if;
	if (ll=23 and cc>=214 and cc<238) then grbp<="010";
	end if;
	if (ll=24 and cc>=27 and cc<168) then grbp<="010";
	end if;
	if (cc=189 and ll=24) then grbp<="010";
	end if;
	if (cc=195 and ll=24) then grbp<="010";
	end if;
	if (ll=24 and cc>=195 and cc<204) then grbp<="010";
	end if;
	if (ll=24 and cc>=214 and cc<237) then grbp<="010";
	end if;
	if (ll=25 and cc>=27 and cc<168) then grbp<="010";
	end if;
	if (cc=194 and ll=25) then grbp<="010";
	end if;
	if (cc=196 and ll=25) then grbp<="010";
	end if;
	if (ll=25 and cc>=196 and cc<204) then grbp<="010";
	end if;
	if (ll=25 and cc>=215 and cc<237) then grbp<="010";
	end if;
	if (ll=26 and cc>=27 and cc<168) then grbp<="010";
	end if;
	if (ll=26 and cc>=198 and cc<205) then grbp<="010";
	end if;
	if (ll=26 and cc>=215 and cc<236) then grbp<="010";
	end if;
	if (ll=27 and cc>=27 and cc<169) then grbp<="010";
	end if;
	if (cc=198 and ll=27) then grbp<="010";
	end if;
	if (ll=27 and cc>=198 and cc<205) then grbp<="010";
	end if;
	if (ll=27 and cc>=216 and cc<235) then grbp<="010";
	end if;
	if (ll=28 and cc>=27 and cc<169) then grbp<="010";
	end if;
	if (ll=28 and cc>=197 and cc<206) then grbp<="010";
	end if;
	if (ll=28 and cc>=216 and cc<235) then grbp<="010";
	end if;
	if (ll=29 and cc>=26 and cc<170) then grbp<="010";
	end if;
	if (cc=191 and ll=29) then grbp<="010";
	end if;
	if (cc=197 and ll=29) then grbp<="010";
	end if;
	if (ll=29 and cc>=197 and cc<206) then grbp<="010";
	end if;
	if (ll=29 and cc>=216 and cc<234) then grbp<="010";
	end if;
	if (ll=30 and cc>=27 and cc<170) then grbp<="010";
	end if;
	if (cc=186 and ll=30) then grbp<="010";
	end if;
	if (cc=191 and ll=30) then grbp<="010";
	end if;
	if (cc=194 and ll=30) then grbp<="010";
	end if;
	if (cc=197 and ll=30) then grbp<="010";
	end if;
	if (ll=30 and cc>=197 and cc<206) then grbp<="010";
	end if;
	if (ll=30 and cc>=217 and cc<234) then grbp<="010";
	end if;
	if (ll=31 and cc>=27 and cc<171) then grbp<="010";
	end if;
	if (cc=194 and ll=31) then grbp<="010";
	end if;
	if (ll=31 and cc>=194 and cc<196) then grbp<="010";
	end if;
	if (ll=31 and cc>=197 and cc<207) then grbp<="010";
	end if;
	if (ll=31 and cc>=217 and cc<233) then grbp<="010";
	end if;
	if (ll=32 and cc>=26 and cc<172) then grbp<="010";
	end if;
	if (ll=32 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (ll=32 and cc>=194 and cc<207) then grbp<="010";
	end if;
	if (ll=32 and cc>=217 and cc<232) then grbp<="010";
	end if;
	if (ll=33 and cc>=27 and cc<171) then grbp<="010";
	end if;
	if (cc=181 and ll=33) then grbp<="010";
	end if;
	if (cc=183 and ll=33) then grbp<="010";
	end if;
	if (cc=186 and ll=33) then grbp<="010";
	end if;
	if (ll=33 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (ll=33 and cc>=195 and cc<207) then grbp<="010";
	end if;
	if (ll=33 and cc>=218 and cc<232) then grbp<="010";
	end if;
	if (ll=34 and cc>=27 and cc<171) then grbp<="010";
	end if;
	if (cc=186 and ll=34) then grbp<="010";
	end if;
	if (ll=34 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (ll=34 and cc>=195 and cc<208) then grbp<="010";
	end if;
	if (ll=34 and cc>=218 and cc<231) then grbp<="010";
	end if;
	if (ll=35 and cc>=27 and cc<174) then grbp<="010";
	end if;
	if (cc=183 and ll=35) then grbp<="010";
	end if;
	if (ll=35 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=35 and cc>=188 and cc<191) then grbp<="010";
	end if;
	if (ll=35 and cc>=194 and cc<208) then grbp<="010";
	end if;
	if (ll=35 and cc>=218 and cc<231) then grbp<="010";
	end if;
	if (ll=36 and cc>=27 and cc<175) then grbp<="010";
	end if;
	if (ll=36 and cc>=179 and cc<181) then grbp<="010";
	end if;
	if (cc=185 and ll=36) then grbp<="010";
	end if;
	if (cc=189 and ll=36) then grbp<="010";
	end if;
	if (ll=36 and cc>=189 and cc<191) then grbp<="010";
	end if;
	if (ll=36 and cc>=193 and cc<208) then grbp<="010";
	end if;
	if (ll=36 and cc>=219 and cc<230) then grbp<="010";
	end if;
	if (cc=27 and ll=37) then grbp<="010";
	end if;
	if (ll=37 and cc>=27 and cc<109) then grbp<="010";
	end if;
	if (cc=112 and ll=37) then grbp<="010";
	end if;
	if (cc=114 and ll=37) then grbp<="010";
	end if;
	if (ll=37 and cc>=114 and cc<175) then grbp<="010";
	end if;
	if (cc=182 and ll=37) then grbp<="010";
	end if;
	if (cc=185 and ll=37) then grbp<="010";
	end if;
	if (cc=188 and ll=37) then grbp<="010";
	end if;
	if (cc=190 and ll=37) then grbp<="010";
	end if;
	if (cc=193 and ll=37) then grbp<="010";
	end if;
	if (ll=37 and cc>=193 and cc<209) then grbp<="010";
	end if;
	if (ll=37 and cc>=219 and cc<230) then grbp<="010";
	end if;
	if (ll=38 and cc>=12 and cc<17) then grbp<="010";
	end if;
	if (ll=38 and cc>=26 and cc<108) then grbp<="010";
	end if;
	if (ll=38 and cc>=118 and cc<175) then grbp<="010";
	end if;
	if (ll=38 and cc>=180 and cc<184) then grbp<="010";
	end if;
	if (cc=190 and ll=38) then grbp<="010";
	end if;
	if (cc=192 and ll=38) then grbp<="010";
	end if;
	if (ll=38 and cc>=192 and cc<209) then grbp<="010";
	end if;
	if (ll=38 and cc>=219 and cc<229) then grbp<="010";
	end if;
	if (ll=39 and cc>=11 and cc<17) then grbp<="010";
	end if;
	if (ll=39 and cc>=27 and cc<102) then grbp<="010";
	end if;
	if (cc=105 and ll=39) then grbp<="010";
	end if;
	if (cc=119 and ll=39) then grbp<="010";
	end if;
	if (ll=39 and cc>=119 and cc<175) then grbp<="010";
	end if;
	if (ll=39 and cc>=180 and cc<183) then grbp<="010";
	end if;
	if (ll=39 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=39 and cc>=187 and cc<189) then grbp<="010";
	end if;
	if (ll=39 and cc>=190 and cc<209) then grbp<="010";
	end if;
	if (ll=39 and cc>=220 and cc<228) then grbp<="010";
	end if;
	if (ll=40 and cc>=11 and cc<17) then grbp<="010";
	end if;
	if (ll=40 and cc>=26 and cc<100) then grbp<="010";
	end if;
	if (ll=40 and cc>=122 and cc<176) then grbp<="010";
	end if;
	if (cc=179 and ll=40) then grbp<="010";
	end if;
	if (cc=181 and ll=40) then grbp<="010";
	end if;
	if (ll=40 and cc>=181 and cc<187) then grbp<="010";
	end if;
	if (cc=190 and ll=40) then grbp<="010";
	end if;
	if (ll=40 and cc>=190 and cc<210) then grbp<="010";
	end if;
	if (ll=40 and cc>=220 and cc<228) then grbp<="010";
	end if;
	if (ll=41 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=41 and cc>=27 and cc<97) then grbp<="010";
	end if;
	if (ll=41 and cc>=123 and cc<177) then grbp<="010";
	end if;
	if (ll=41 and cc>=178 and cc<186) then grbp<="010";
	end if;
	if (cc=190 and ll=41) then grbp<="010";
	end if;
	if (ll=41 and cc>=190 and cc<210) then grbp<="010";
	end if;
	if (ll=41 and cc>=220 and cc<227) then grbp<="010";
	end if;
	if (ll=42 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=42 and cc>=27 and cc<95) then grbp<="010";
	end if;
	if (ll=42 and cc>=125 and cc<177) then grbp<="010";
	end if;
	if (cc=180 and ll=42) then grbp<="010";
	end if;
	if (cc=183 and ll=42) then grbp<="010";
	end if;
	if (ll=42 and cc>=183 and cc<189) then grbp<="010";
	end if;
	if (ll=42 and cc>=190 and cc<210) then grbp<="010";
	end if;
	if (ll=42 and cc>=221 and cc<227) then grbp<="010";
	end if;
	if (ll=43 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=43 and cc>=27 and cc<93) then grbp<="010";
	end if;
	if (cc=127 and ll=43) then grbp<="010";
	end if;
	if (ll=43 and cc>=127 and cc<178) then grbp<="010";
	end if;
	if (ll=43 and cc>=180 and cc<184) then grbp<="010";
	end if;
	if (ll=43 and cc>=185 and cc<211) then grbp<="010";
	end if;
	if (ll=43 and cc>=221 and cc<226) then grbp<="010";
	end if;
	if (ll=44 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=44 and cc>=27 and cc<96) then grbp<="010";
	end if;
	if (ll=44 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=44 and cc>=128 and cc<211) then grbp<="010";
	end if;
	if (ll=44 and cc>=221 and cc<225) then grbp<="010";
	end if;
	if (ll=45 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=45 and cc>=27 and cc<93) then grbp<="010";
	end if;
	if (cc=99 and ll=45) then grbp<="010";
	end if;
	if (ll=45 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (ll=45 and cc>=129 and cc<179) then grbp<="010";
	end if;
	if (ll=45 and cc>=180 and cc<212) then grbp<="010";
	end if;
	if (ll=45 and cc>=222 and cc<225) then grbp<="010";
	end if;
	if (ll=46 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=46 and cc>=27 and cc<92) then grbp<="010";
	end if;
	if (cc=97 and ll=46) then grbp<="010";
	end if;
	if (cc=100 and ll=46) then grbp<="010";
	end if;
	if (cc=102 and ll=46) then grbp<="010";
	end if;
	if (cc=130 and ll=46) then grbp<="010";
	end if;
	if (ll=46 and cc>=130 and cc<212) then grbp<="010";
	end if;
	if (ll=46 and cc>=222 and cc<224) then grbp<="010";
	end if;
	if (ll=47 and cc>=8 and cc<17) then grbp<="010";
	end if;
	if (ll=47 and cc>=27 and cc<86) then grbp<="010";
	end if;
	if (ll=47 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (cc=95 and ll=47) then grbp<="010";
	end if;
	if (cc=97 and ll=47) then grbp<="010";
	end if;
	if (ll=47 and cc>=97 and cc<100) then grbp<="010";
	end if;
	if (ll=47 and cc>=131 and cc<181) then grbp<="010";
	end if;
	if (ll=47 and cc>=182 and cc<212) then grbp<="010";
	end if;
	if (ll=47 and cc>=222 and cc<224) then grbp<="010";
	end if;
	if (ll=48 and cc>=8 and cc<17) then grbp<="010";
	end if;
	if (ll=48 and cc>=27 and cc<83) then grbp<="010";
	end if;
	if (ll=48 and cc>=87 and cc<95) then grbp<="010";
	end if;
	if (ll=48 and cc>=96 and cc<99) then grbp<="010";
	end if;
	if (cc=132 and ll=48) then grbp<="010";
	end if;
	if (ll=48 and cc>=132 and cc<181) then grbp<="010";
	end if;
	if (ll=48 and cc>=182 and cc<213) then grbp<="010";
	end if;
	if (cc=7 and ll=49) then grbp<="010";
	end if;
	if (ll=49 and cc>=7 and cc<16) then grbp<="010";
	end if;
	if (ll=49 and cc>=27 and cc<81) then grbp<="010";
	end if;
	if (cc=86 and ll=49) then grbp<="010";
	end if;
	if (ll=49 and cc>=86 and cc<99) then grbp<="010";
	end if;
	if (cc=132 and ll=49) then grbp<="010";
	end if;
	if (ll=49 and cc>=132 and cc<179) then grbp<="010";
	end if;
	if (ll=49 and cc>=180 and cc<213) then grbp<="010";
	end if;
	if (ll=50 and cc>=7 and cc<16) then grbp<="010";
	end if;
	if (ll=50 and cc>=27 and cc<80) then grbp<="010";
	end if;
	if (ll=50 and cc>=84 and cc<101) then grbp<="010";
	end if;
	if (cc=133 and ll=50) then grbp<="010";
	end if;
	if (ll=50 and cc>=133 and cc<213) then grbp<="010";
	end if;
	if (ll=51 and cc>=7 and cc<17) then grbp<="010";
	end if;
	if (ll=51 and cc>=27 and cc<101) then grbp<="010";
	end if;
	if (cc=134 and ll=51) then grbp<="010";
	end if;
	if (ll=51 and cc>=134 and cc<214) then grbp<="010";
	end if;
	if (cc=7 and ll=52) then grbp<="010";
	end if;
	if (ll=52 and cc>=7 and cc<16) then grbp<="010";
	end if;
	if (ll=52 and cc>=27 and cc<78) then grbp<="010";
	end if;
	if (ll=52 and cc>=79 and cc<103) then grbp<="010";
	end if;
	if (ll=52 and cc>=135 and cc<183) then grbp<="010";
	end if;
	if (ll=52 and cc>=184 and cc<214) then grbp<="010";
	end if;
	if (cc=7 and ll=53) then grbp<="010";
	end if;
	if (ll=53 and cc>=7 and cc<16) then grbp<="010";
	end if;
	if (ll=53 and cc>=27 and cc<77) then grbp<="010";
	end if;
	if (ll=53 and cc>=79 and cc<102) then grbp<="010";
	end if;
	if (cc=136 and ll=53) then grbp<="010";
	end if;
	if (ll=53 and cc>=136 and cc<214) then grbp<="010";
	end if;
	if (ll=54 and cc>=6 and cc<16) then grbp<="010";
	end if;
	if (ll=54 and cc>=27 and cc<77) then grbp<="010";
	end if;
	if (ll=54 and cc>=78 and cc<103) then grbp<="010";
	end if;
	if (cc=137 and ll=54) then grbp<="010";
	end if;
	if (ll=54 and cc>=137 and cc<215) then grbp<="010";
	end if;
	if (cc=6 and ll=55) then grbp<="010";
	end if;
	if (ll=55 and cc>=6 and cc<16) then grbp<="010";
	end if;
	if (ll=55 and cc>=27 and cc<77) then grbp<="010";
	end if;
	if (ll=55 and cc>=78 and cc<102) then grbp<="010";
	end if;
	if (cc=137 and ll=55) then grbp<="010";
	end if;
	if (ll=55 and cc>=137 and cc<215) then grbp<="010";
	end if;
	if (ll=56 and cc>=5 and cc<16) then grbp<="010";
	end if;
	if (ll=56 and cc>=26 and cc<77) then grbp<="010";
	end if;
	if (ll=56 and cc>=78 and cc<104) then grbp<="010";
	end if;
	if (ll=56 and cc>=105 and cc<107) then grbp<="010";
	end if;
	if (ll=56 and cc>=138 and cc<215) then grbp<="010";
	end if;
	if (cc=5 and ll=57) then grbp<="010";
	end if;
	if (ll=57 and cc>=5 and cc<16) then grbp<="010";
	end if;
	if (ll=57 and cc>=26 and cc<106) then grbp<="010";
	end if;
	if (ll=57 and cc>=139 and cc<216) then grbp<="010";
	end if;
	if (cc=5 and ll=58) then grbp<="010";
	end if;
	if (ll=58 and cc>=5 and cc<17) then grbp<="010";
	end if;
	if (ll=58 and cc>=26 and cc<105) then grbp<="010";
	end if;
	if (cc=140 and ll=58) then grbp<="010";
	end if;
	if (ll=58 and cc>=140 and cc<216) then grbp<="010";
	end if;
	if (cc=5 and ll=59) then grbp<="010";
	end if;
	if (ll=59 and cc>=5 and cc<17) then grbp<="010";
	end if;
	if (ll=59 and cc>=26 and cc<106) then grbp<="010";
	end if;
	if (cc=141 and ll=59) then grbp<="010";
	end if;
	if (ll=59 and cc>=141 and cc<214) then grbp<="010";
	end if;
	if (cc=218 and ll=59) then grbp<="010";
	end if;
	if (cc=4 and ll=60) then grbp<="010";
	end if;
	if (ll=60 and cc>=4 and cc<17) then grbp<="010";
	end if;
	if (ll=60 and cc>=26 and cc<108) then grbp<="010";
	end if;
	if (ll=60 and cc>=141 and cc<214) then grbp<="010";
	end if;
	if (cc=250 and ll=60) then grbp<="010";
	end if;
	if (cc=4 and ll=61) then grbp<="010";
	end if;
	if (ll=61 and cc>=4 and cc<17) then grbp<="010";
	end if;
	if (ll=61 and cc>=26 and cc<107) then grbp<="010";
	end if;
	if (cc=142 and ll=61) then grbp<="010";
	end if;
	if (ll=61 and cc>=142 and cc<214) then grbp<="010";
	end if;
	if (ll=61 and cc>=215 and cc<218) then grbp<="010";
	end if;
	if (cc=4 and ll=62) then grbp<="010";
	end if;
	if (ll=62 and cc>=4 and cc<16) then grbp<="010";
	end if;
	if (ll=62 and cc>=26 and cc<74) then grbp<="010";
	end if;
	if (ll=62 and cc>=75 and cc<106) then grbp<="010";
	end if;
	if (cc=144 and ll=62) then grbp<="010";
	end if;
	if (ll=62 and cc>=144 and cc<170) then grbp<="010";
	end if;
	if (ll=62 and cc>=172 and cc<217) then grbp<="010";
	end if;
	if (ll=62 and cc>=249 and cc<251) then grbp<="010";
	end if;
	if (cc=3 and ll=63) then grbp<="010";
	end if;
	if (ll=63 and cc>=3 and cc<17) then grbp<="010";
	end if;
	if (ll=63 and cc>=26 and cc<74) then grbp<="010";
	end if;
	if (ll=63 and cc>=75 and cc<106) then grbp<="010";
	end if;
	if (cc=109 and ll=63) then grbp<="010";
	end if;
	if (cc=145 and ll=63) then grbp<="010";
	end if;
	if (ll=63 and cc>=145 and cc<168) then grbp<="010";
	end if;
	if (ll=63 and cc>=170 and cc<213) then grbp<="010";
	end if;
	if (ll=63 and cc>=215 and cc<217) then grbp<="010";
	end if;
	if (cc=3 and ll=64) then grbp<="010";
	end if;
	if (ll=64 and cc>=3 and cc<16) then grbp<="010";
	end if;
	if (ll=64 and cc>=27 and cc<74) then grbp<="010";
	end if;
	if (ll=64 and cc>=75 and cc<105) then grbp<="010";
	end if;
	if (ll=64 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=64 and cc>=146 and cc<168) then grbp<="010";
	end if;
	if (cc=171 and ll=64) then grbp<="010";
	end if;
	if (ll=64 and cc>=171 and cc<213) then grbp<="010";
	end if;
	if (ll=64 and cc>=215 and cc<217) then grbp<="010";
	end if;
	if (ll=64 and cc>=248 and cc<250) then grbp<="010";
	end if;
	if (ll=65 and cc>=2 and cc<16) then grbp<="010";
	end if;
	if (ll=65 and cc>=27 and cc<108) then grbp<="010";
	end if;
	if (cc=146 and ll=65) then grbp<="010";
	end if;
	if (ll=65 and cc>=146 and cc<168) then grbp<="010";
	end if;
	if (ll=65 and cc>=169 and cc<212) then grbp<="010";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="010";
	end if;
	if (ll=65 and cc>=248 and cc<250) then grbp<="010";
	end if;
	if (ll=66 and cc>=2 and cc<16) then grbp<="010";
	end if;
	if (ll=66 and cc>=26 and cc<105) then grbp<="010";
	end if;
	if (ll=66 and cc>=106 and cc<108) then grbp<="010";
	end if;
	if (cc=146 and ll=66) then grbp<="010";
	end if;
	if (ll=66 and cc>=146 and cc<169) then grbp<="010";
	end if;
	if (ll=66 and cc>=170 and cc<212) then grbp<="010";
	end if;
	if (ll=66 and cc>=213 and cc<216) then grbp<="010";
	end if;
	if (ll=66 and cc>=247 and cc<249) then grbp<="010";
	end if;
	if (ll=67 and cc>=2 and cc<17) then grbp<="010";
	end if;
	if (ll=67 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (cc=147 and ll=67) then grbp<="010";
	end if;
	if (ll=67 and cc>=147 and cc<215) then grbp<="010";
	end if;
	if (ll=67 and cc>=247 and cc<249) then grbp<="010";
	end if;
	if (ll=68 and cc>=2 and cc<16) then grbp<="010";
	end if;
	if (ll=68 and cc>=27 and cc<109) then grbp<="010";
	end if;
	if (ll=68 and cc>=147 and cc<211) then grbp<="010";
	end if;
	if (ll=68 and cc>=213 and cc<215) then grbp<="010";
	end if;
	if (ll=68 and cc>=246 and cc<249) then grbp<="010";
	end if;
	if (ll=69 and cc>=1 and cc<17) then grbp<="010";
	end if;
	if (ll=69 and cc>=26 and cc<108) then grbp<="010";
	end if;
	if (cc=148 and ll=69) then grbp<="010";
	end if;
	if (ll=69 and cc>=148 and cc<169) then grbp<="010";
	end if;
	if (ll=69 and cc>=170 and cc<214) then grbp<="010";
	end if;
	if (ll=69 and cc>=246 and cc<249) then grbp<="010";
	end if;
	if (ll=70 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=70 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (ll=70 and cc>=148 and cc<168) then grbp<="010";
	end if;
	if (ll=70 and cc>=169 and cc<214) then grbp<="010";
	end if;
	if (ll=70 and cc>=245 and cc<250) then grbp<="010";
	end if;
	if (ll=71 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=71 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (cc=148 and ll=71) then grbp<="010";
	end if;
	if (ll=71 and cc>=148 and cc<168) then grbp<="010";
	end if;
	if (ll=71 and cc>=169 and cc<181) then grbp<="010";
	end if;
	if (ll=71 and cc>=183 and cc<214) then grbp<="010";
	end if;
	if (ll=71 and cc>=244 and cc<247) then grbp<="010";
	end if;
	if (ll=71 and cc>=248 and cc<250) then grbp<="010";
	end if;
	if (ll=72 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=72 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (ll=72 and cc>=149 and cc<181) then grbp<="010";
	end if;
	if (ll=72 and cc>=183 and cc<213) then grbp<="010";
	end if;
	if (ll=72 and cc>=244 and cc<247) then grbp<="010";
	end if;
	if (ll=72 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=73) then grbp<="010";
	end if;
	if (ll=73 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=73 and cc>=26 and cc<107) then grbp<="010";
	end if;
	if (ll=73 and cc>=149 and cc<168) then grbp<="010";
	end if;
	if (ll=73 and cc>=169 and cc<181) then grbp<="010";
	end if;
	if (ll=73 and cc>=183 and cc<213) then grbp<="010";
	end if;
	if (ll=73 and cc>=243 and cc<246) then grbp<="010";
	end if;
	if (ll=73 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=74) then grbp<="010";
	end if;
	if (ll=74 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=74 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (ll=74 and cc>=150 and cc<181) then grbp<="010";
	end if;
	if (ll=74 and cc>=184 and cc<212) then grbp<="010";
	end if;
	if (ll=74 and cc>=242 and cc<246) then grbp<="010";
	end if;
	if (ll=74 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=75) then grbp<="010";
	end if;
	if (ll=75 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=75 and cc>=26 and cc<110) then grbp<="010";
	end if;
	if (ll=75 and cc>=150 and cc<170) then grbp<="010";
	end if;
	if (ll=75 and cc>=171 and cc<181) then grbp<="010";
	end if;
	if (ll=75 and cc>=184 and cc<212) then grbp<="010";
	end if;
	if (ll=75 and cc>=242 and cc<246) then grbp<="010";
	end if;
	if (ll=75 and cc>=248 and cc<250) then grbp<="010";
	end if;
	if (ll=76 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=76 and cc>=27 and cc<111) then grbp<="010";
	end if;
	if (ll=76 and cc>=151 and cc<168) then grbp<="010";
	end if;
	if (ll=76 and cc>=169 and cc<181) then grbp<="010";
	end if;
	if (ll=76 and cc>=184 and cc<212) then grbp<="010";
	end if;
	if (ll=76 and cc>=241 and cc<245) then grbp<="010";
	end if;
	if (ll=76 and cc>=248 and cc<250) then grbp<="010";
	end if;
	if (ll=77 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=77 and cc>=26 and cc<111) then grbp<="010";
	end if;
	if (ll=77 and cc>=151 and cc<181) then grbp<="010";
	end if;
	if (ll=77 and cc>=185 and cc<211) then grbp<="010";
	end if;
	if (ll=77 and cc>=240 and cc<246) then grbp<="010";
	end if;
	if (ll=77 and cc>=247 and cc<249) then grbp<="010";
	end if;
	if (ll=78 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=78 and cc>=27 and cc<111) then grbp<="010";
	end if;
	if (ll=78 and cc>=151 and cc<181) then grbp<="010";
	end if;
	if (ll=78 and cc>=185 and cc<211) then grbp<="010";
	end if;
	if (ll=78 and cc>=240 and cc<244) then grbp<="010";
	end if;
	if (ll=78 and cc>=245 and cc<249) then grbp<="010";
	end if;
	if (ll=79 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=79 and cc>=27 and cc<110) then grbp<="010";
	end if;
	if (cc=152 and ll=79) then grbp<="010";
	end if;
	if (ll=79 and cc>=152 and cc<181) then grbp<="010";
	end if;
	if (ll=79 and cc>=185 and cc<210) then grbp<="010";
	end if;
	if (ll=79 and cc>=240 and cc<244) then grbp<="010";
	end if;
	if (ll=79 and cc>=245 and cc<248) then grbp<="010";
	end if;
	if (ll=80 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=80 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (cc=153 and ll=80) then grbp<="010";
	end if;
	if (ll=80 and cc>=153 and cc<181) then grbp<="010";
	end if;
	if (ll=80 and cc>=186 and cc<210) then grbp<="010";
	end if;
	if (ll=80 and cc>=239 and cc<248) then grbp<="010";
	end if;
	if (ll=81 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=81 and cc>=26 and cc<109) then grbp<="010";
	end if;
	if (cc=114 and ll=81) then grbp<="010";
	end if;
	if (ll=81 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (ll=81 and cc>=154 and cc<168) then grbp<="010";
	end if;
	if (ll=81 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (ll=81 and cc>=172 and cc<181) then grbp<="010";
	end if;
	if (ll=81 and cc>=186 and cc<210) then grbp<="010";
	end if;
	if (ll=81 and cc>=239 and cc<244) then grbp<="010";
	end if;
	if (ll=81 and cc>=245 and cc<247) then grbp<="010";
	end if;
	if (ll=82 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=82 and cc>=26 and cc<111) then grbp<="010";
	end if;
	if (cc=155 and ll=82) then grbp<="010";
	end if;
	if (ll=82 and cc>=155 and cc<175) then grbp<="010";
	end if;
	if (ll=82 and cc>=176 and cc<181) then grbp<="010";
	end if;
	if (ll=82 and cc>=187 and cc<209) then grbp<="010";
	end if;
	if (ll=82 and cc>=239 and cc<242) then grbp<="010";
	end if;
	if (cc=245 and ll=82) then grbp<="010";
	end if;
	if (ll=82 and cc>=245 and cc<247) then grbp<="010";
	end if;
	if (ll=83 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=83 and cc>=26 and cc<110) then grbp<="010";
	end if;
	if (cc=155 and ll=83) then grbp<="010";
	end if;
	if (ll=83 and cc>=155 and cc<168) then grbp<="010";
	end if;
	if (ll=83 and cc>=169 and cc<175) then grbp<="010";
	end if;
	if (ll=83 and cc>=176 and cc<181) then grbp<="010";
	end if;
	if (ll=83 and cc>=187 and cc<209) then grbp<="010";
	end if;
	if (ll=83 and cc>=238 and cc<243) then grbp<="010";
	end if;
	if (ll=83 and cc>=244 and cc<246) then grbp<="010";
	end if;
	if (ll=84 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=84 and cc>=26 and cc<111) then grbp<="010";
	end if;
	if (cc=156 and ll=84) then grbp<="010";
	end if;
	if (cc=158 and ll=84) then grbp<="010";
	end if;
	if (ll=84 and cc>=158 and cc<181) then grbp<="010";
	end if;
	if (ll=84 and cc>=187 and cc<209) then grbp<="010";
	end if;
	if (ll=84 and cc>=237 and cc<246) then grbp<="010";
	end if;
	if (ll=85 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=85 and cc>=26 and cc<113) then grbp<="010";
	end if;
	if (cc=158 and ll=85) then grbp<="010";
	end if;
	if (ll=85 and cc>=158 and cc<168) then grbp<="010";
	end if;
	if (ll=85 and cc>=169 and cc<181) then grbp<="010";
	end if;
	if (ll=85 and cc>=187 and cc<208) then grbp<="010";
	end if;
	if (ll=85 and cc>=237 and cc<239) then grbp<="010";
	end if;
	if (ll=85 and cc>=240 and cc<245) then grbp<="010";
	end if;
	if (ll=86 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=86 and cc>=27 and cc<112) then grbp<="010";
	end if;
	if (ll=86 and cc>=159 and cc<181) then grbp<="010";
	end if;
	if (ll=86 and cc>=188 and cc<208) then grbp<="010";
	end if;
	if (ll=86 and cc>=236 and cc<245) then grbp<="010";
	end if;
	if (ll=87 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=87 and cc>=26 and cc<111) then grbp<="010";
	end if;
	if (cc=159 and ll=87) then grbp<="010";
	end if;
	if (ll=87 and cc>=159 and cc<181) then grbp<="010";
	end if;
	if (ll=87 and cc>=188 and cc<207) then grbp<="010";
	end if;
	if (ll=87 and cc>=236 and cc<239) then grbp<="010";
	end if;
	if (ll=87 and cc>=240 and cc<244) then grbp<="010";
	end if;
	if (ll=88 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=88 and cc>=27 and cc<64) then grbp<="010";
	end if;
	if (ll=88 and cc>=65 and cc<110) then grbp<="010";
	end if;
	if (ll=88 and cc>=160 and cc<181) then grbp<="010";
	end if;
	if (ll=88 and cc>=189 and cc<207) then grbp<="010";
	end if;
	if (ll=88 and cc>=236 and cc<238) then grbp<="010";
	end if;
	if (ll=88 and cc>=240 and cc<243) then grbp<="010";
	end if;
	if (ll=89 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=89 and cc>=27 and cc<64) then grbp<="010";
	end if;
	if (ll=89 and cc>=65 and cc<109) then grbp<="010";
	end if;
	if (ll=89 and cc>=159 and cc<181) then grbp<="010";
	end if;
	if (ll=89 and cc>=189 and cc<207) then grbp<="010";
	end if;
	if (ll=89 and cc>=235 and cc<238) then grbp<="010";
	end if;
	if (ll=89 and cc>=239 and cc<243) then grbp<="010";
	end if;
	if (ll=90 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=90 and cc>=27 and cc<64) then grbp<="010";
	end if;
	if (ll=90 and cc>=65 and cc<108) then grbp<="010";
	end if;
	if (ll=90 and cc>=158 and cc<171) then grbp<="010";
	end if;
	if (ll=90 and cc>=172 and cc<181) then grbp<="010";
	end if;
	if (ll=90 and cc>=190 and cc<206) then grbp<="010";
	end if;
	if (ll=90 and cc>=235 and cc<243) then grbp<="010";
	end if;
	if (ll=91 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=91 and cc>=27 and cc<64) then grbp<="010";
	end if;
	if (ll=91 and cc>=65 and cc<108) then grbp<="010";
	end if;
	if (cc=161 and ll=91) then grbp<="010";
	end if;
	if (ll=91 and cc>=161 and cc<172) then grbp<="010";
	end if;
	if (ll=91 and cc>=173 and cc<181) then grbp<="010";
	end if;
	if (ll=91 and cc>=190 and cc<206) then grbp<="010";
	end if;
	if (ll=91 and cc>=234 and cc<242) then grbp<="010";
	end if;
	if (ll=92 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=92 and cc>=27 and cc<63) then grbp<="010";
	end if;
	if (ll=92 and cc>=65 and cc<107) then grbp<="010";
	end if;
	if (cc=161 and ll=92) then grbp<="010";
	end if;
	if (ll=92 and cc>=161 and cc<181) then grbp<="010";
	end if;
	if (ll=92 and cc>=191 and cc<194) then grbp<="010";
	end if;
	if (ll=92 and cc>=199 and cc<201) then grbp<="010";
	end if;
	if (ll=92 and cc>=202 and cc<205) then grbp<="010";
	end if;
	if (cc=237 and ll=92) then grbp<="010";
	end if;
	if (ll=92 and cc>=237 and cc<242) then grbp<="010";
	end if;
	if (ll=93 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=93 and cc>=27 and cc<63) then grbp<="010";
	end if;
	if (ll=93 and cc>=65 and cc<106) then grbp<="010";
	end if;
	if (ll=93 and cc>=161 and cc<174) then grbp<="010";
	end if;
	if (ll=93 and cc>=176 and cc<181) then grbp<="010";
	end if;
	if (ll=93 and cc>=191 and cc<193) then grbp<="010";
	end if;
	if (ll=93 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (ll=93 and cc>=234 and cc<242) then grbp<="010";
	end if;
	if (ll=94 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=94 and cc>=27 and cc<63) then grbp<="010";
	end if;
	if (ll=94 and cc>=65 and cc<106) then grbp<="010";
	end if;
	if (ll=94 and cc>=161 and cc<181) then grbp<="010";
	end if;
	if (ll=94 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (ll=94 and cc>=233 and cc<241) then grbp<="010";
	end if;
	if (ll=95 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=95 and cc>=27 and cc<63) then grbp<="010";
	end if;
	if (ll=95 and cc>=65 and cc<104) then grbp<="010";
	end if;
	if (ll=95 and cc>=162 and cc<181) then grbp<="010";
	end if;
	if (cc=233 and ll=95) then grbp<="010";
	end if;
	if (ll=95 and cc>=233 and cc<235) then grbp<="010";
	end if;
	if (ll=95 and cc>=236 and cc<241) then grbp<="010";
	end if;
	if (ll=96 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=96 and cc>=26 and cc<62) then grbp<="010";
	end if;
	if (ll=96 and cc>=65 and cc<104) then grbp<="010";
	end if;
	if (cc=162 and ll=96) then grbp<="010";
	end if;
	if (ll=96 and cc>=162 and cc<181) then grbp<="010";
	end if;
	if (ll=96 and cc>=232 and cc<240) then grbp<="010";
	end if;
	if (ll=97 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=97 and cc>=26 and cc<62) then grbp<="010";
	end if;
	if (ll=97 and cc>=64 and cc<103) then grbp<="010";
	end if;
	if (cc=162 and ll=97) then grbp<="010";
	end if;
	if (ll=97 and cc>=162 and cc<181) then grbp<="010";
	end if;
	if (cc=234 and ll=97) then grbp<="010";
	end if;
	if (cc=236 and ll=97) then grbp<="010";
	end if;
	if (ll=97 and cc>=236 and cc<239) then grbp<="010";
	end if;
	if (ll=98 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=98 and cc>=27 and cc<62) then grbp<="010";
	end if;
	if (ll=98 and cc>=64 and cc<102) then grbp<="010";
	end if;
	if (ll=98 and cc>=162 and cc<181) then grbp<="010";
	end if;
	if (ll=98 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=98 and cc>=234 and cc<239) then grbp<="010";
	end if;
	if (ll=99 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=99 and cc>=27 and cc<62) then grbp<="010";
	end if;
	if (ll=99 and cc>=64 and cc<101) then grbp<="010";
	end if;
	if (ll=99 and cc>=161 and cc<181) then grbp<="010";
	end if;
	if (cc=235 and ll=99) then grbp<="010";
	end if;
	if (ll=99 and cc>=235 and cc<238) then grbp<="010";
	end if;
	if (ll=100 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=100 and cc>=27 and cc<62) then grbp<="010";
	end if;
	if (ll=100 and cc>=65 and cc<101) then grbp<="010";
	end if;
	if (ll=100 and cc>=161 and cc<172) then grbp<="010";
	end if;
	if (ll=100 and cc>=173 and cc<181) then grbp<="010";
	end if;
	if (ll=100 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=100 and cc>=234 and cc<238) then grbp<="010";
	end if;
	if (ll=101 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=101 and cc>=27 and cc<61) then grbp<="010";
	end if;
	if (ll=101 and cc>=64 and cc<100) then grbp<="010";
	end if;
	if (ll=101 and cc>=162 and cc<168) then grbp<="010";
	end if;
	if (cc=171 and ll=101) then grbp<="010";
	end if;
	if (ll=101 and cc>=171 and cc<181) then grbp<="010";
	end if;
	if (cc=232 and ll=101) then grbp<="010";
	end if;
	if (cc=234 and ll=101) then grbp<="010";
	end if;
	if (ll=101 and cc>=234 and cc<238) then grbp<="010";
	end if;
	if (ll=102 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=102 and cc>=27 and cc<61) then grbp<="010";
	end if;
	if (ll=102 and cc>=64 and cc<99) then grbp<="010";
	end if;
	if (ll=102 and cc>=162 and cc<168) then grbp<="010";
	end if;
	if (ll=102 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (ll=102 and cc>=172 and cc<181) then grbp<="010";
	end if;
	if (cc=233 and ll=102) then grbp<="010";
	end if;
	if (ll=102 and cc>=233 and cc<237) then grbp<="010";
	end if;
	if (ll=103 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=103 and cc>=26 and cc<61) then grbp<="010";
	end if;
	if (ll=103 and cc>=64 and cc<98) then grbp<="010";
	end if;
	if (ll=103 and cc>=163 and cc<168) then grbp<="010";
	end if;
	if (cc=175 and ll=103) then grbp<="010";
	end if;
	if (ll=103 and cc>=175 and cc<181) then grbp<="010";
	end if;
	if (ll=103 and cc>=229 and cc<231) then grbp<="010";
	end if;
	if (ll=103 and cc>=233 and cc<237) then grbp<="010";
	end if;
	if (ll=104 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=104 and cc>=27 and cc<61) then grbp<="010";
	end if;
	if (ll=104 and cc>=64 and cc<98) then grbp<="010";
	end if;
	if (ll=104 and cc>=163 and cc<171) then grbp<="010";
	end if;
	if (cc=175 and ll=104) then grbp<="010";
	end if;
	if (ll=104 and cc>=175 and cc<181) then grbp<="010";
	end if;
	if (ll=104 and cc>=229 and cc<231) then grbp<="010";
	end if;
	if (ll=104 and cc>=232 and cc<236) then grbp<="010";
	end if;
	if (ll=105 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=105 and cc>=26 and cc<61) then grbp<="010";
	end if;
	if (ll=105 and cc>=64 and cc<97) then grbp<="010";
	end if;
	if (ll=105 and cc>=163 and cc<171) then grbp<="010";
	end if;
	if (ll=105 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=105 and cc>=175 and cc<180) then grbp<="010";
	end if;
	if (cc=232 and ll=105) then grbp<="010";
	end if;
	if (ll=105 and cc>=232 and cc<236) then grbp<="010";
	end if;
	if (ll=106 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=106 and cc>=27 and cc<61) then grbp<="010";
	end if;
	if (ll=106 and cc>=64 and cc<97) then grbp<="010";
	end if;
	if (ll=106 and cc>=164 and cc<169) then grbp<="010";
	end if;
	if (cc=172 and ll=106) then grbp<="010";
	end if;
	if (cc=174 and ll=106) then grbp<="010";
	end if;
	if (ll=106 and cc>=174 and cc<180) then grbp<="010";
	end if;
	if (ll=106 and cc>=228 and cc<230) then grbp<="010";
	end if;
	if (ll=106 and cc>=232 and cc<235) then grbp<="010";
	end if;
	if (ll=107 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=107 and cc>=27 and cc<61) then grbp<="010";
	end if;
	if (ll=107 and cc>=64 and cc<96) then grbp<="010";
	end if;
	if (ll=107 and cc>=164 and cc<171) then grbp<="010";
	end if;
	if (ll=107 and cc>=172 and cc<180) then grbp<="010";
	end if;
	if (ll=107 and cc>=228 and cc<230) then grbp<="010";
	end if;
	if (ll=107 and cc>=232 and cc<235) then grbp<="010";
	end if;
	if (ll=108 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=108 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=108 and cc>=64 and cc<96) then grbp<="010";
	end if;
	if (ll=108 and cc>=165 and cc<171) then grbp<="010";
	end if;
	if (ll=108 and cc>=172 and cc<180) then grbp<="010";
	end if;
	if (cc=228 and ll=108) then grbp<="010";
	end if;
	if (cc=231 and ll=108) then grbp<="010";
	end if;
	if (ll=108 and cc>=231 and cc<234) then grbp<="010";
	end if;
	if (ll=109 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=109 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=109 and cc>=63 and cc<95) then grbp<="010";
	end if;
	if (cc=100 and ll=109) then grbp<="010";
	end if;
	if (cc=105 and ll=109) then grbp<="010";
	end if;
	if (cc=166 and ll=109) then grbp<="010";
	end if;
	if (ll=109 and cc>=166 and cc<172) then grbp<="010";
	end if;
	if (ll=109 and cc>=173 and cc<181) then grbp<="010";
	end if;
	if (ll=109 and cc>=227 and cc<229) then grbp<="010";
	end if;
	if (cc=0 and ll=110) then grbp<="010";
	end if;
	if (ll=110 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=110 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=110 and cc>=63 and cc<94) then grbp<="010";
	end if;
	if (cc=104 and ll=110) then grbp<="010";
	end if;
	if (cc=166 and ll=110) then grbp<="010";
	end if;
	if (ll=110 and cc>=166 and cc<180) then grbp<="010";
	end if;
	if (ll=110 and cc>=227 and cc<229) then grbp<="010";
	end if;
	if (ll=110 and cc>=230 and cc<234) then grbp<="010";
	end if;
	if (ll=111 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=111 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=111 and cc>=63 and cc<94) then grbp<="010";
	end if;
	if (cc=100 and ll=111) then grbp<="010";
	end if;
	if (cc=167 and ll=111) then grbp<="010";
	end if;
	if (ll=111 and cc>=167 and cc<179) then grbp<="010";
	end if;
	if (cc=230 and ll=111) then grbp<="010";
	end if;
	if (cc=232 and ll=111) then grbp<="010";
	end if;
	if (cc=0 and ll=112) then grbp<="010";
	end if;
	if (ll=112 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=112 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=112 and cc>=63 and cc<93) then grbp<="010";
	end if;
	if (ll=112 and cc>=97 and cc<99) then grbp<="010";
	end if;
	if (cc=102 and ll=112) then grbp<="010";
	end if;
	if (cc=167 and ll=112) then grbp<="010";
	end if;
	if (ll=112 and cc>=167 and cc<169) then grbp<="010";
	end if;
	if (ll=112 and cc>=170 and cc<177) then grbp<="010";
	end if;
	if (ll=112 and cc>=226 and cc<228) then grbp<="010";
	end if;
	if (ll=112 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=113 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=113 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=113 and cc>=63 and cc<93) then grbp<="010";
	end if;
	if (ll=113 and cc>=97 and cc<100) then grbp<="010";
	end if;
	if (ll=113 and cc>=101 and cc<103) then grbp<="010";
	end if;
	if (ll=113 and cc>=167 and cc<176) then grbp<="010";
	end if;
	if (ll=113 and cc>=226 and cc<228) then grbp<="010";
	end if;
	if (ll=113 and cc>=229 and cc<232) then grbp<="010";
	end if;
	if (ll=114 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=114 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=114 and cc>=63 and cc<92) then grbp<="010";
	end if;
	if (ll=114 and cc>=95 and cc<100) then grbp<="010";
	end if;
	if (ll=114 and cc>=101 and cc<103) then grbp<="010";
	end if;
	if (ll=114 and cc>=168 and cc<175) then grbp<="010";
	end if;
	if (ll=114 and cc>=225 and cc<228) then grbp<="010";
	end if;
	if (ll=114 and cc>=229 and cc<232) then grbp<="010";
	end if;
	if (ll=115 and cc>=0 and cc<18) then grbp<="010";
	end if;
	if (ll=115 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=115 and cc>=63 and cc<93) then grbp<="010";
	end if;
	if (ll=115 and cc>=95 and cc<98) then grbp<="010";
	end if;
	if (ll=115 and cc>=100 and cc<102) then grbp<="010";
	end if;
	if (ll=115 and cc>=168 and cc<174) then grbp<="010";
	end if;
	if (ll=115 and cc>=225 and cc<227) then grbp<="010";
	end if;
	if (ll=115 and cc>=229 and cc<232) then grbp<="010";
	end if;
	if (ll=116 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=116 and cc>=27 and cc<60) then grbp<="010";
	end if;
	if (ll=116 and cc>=62 and cc<93) then grbp<="010";
	end if;
	if (ll=116 and cc>=95 and cc<98) then grbp<="010";
	end if;
	if (ll=116 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (ll=116 and cc>=168 and cc<173) then grbp<="010";
	end if;
	if (cc=224 and ll=116) then grbp<="010";
	end if;
	if (ll=116 and cc>=224 and cc<227) then grbp<="010";
	end if;
	if (ll=116 and cc>=228 and cc<232) then grbp<="010";
	end if;
	if (ll=117 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=117 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=117 and cc>=63 and cc<89) then grbp<="010";
	end if;
	if (cc=92 and ll=117) then grbp<="010";
	end if;
	if (cc=94 and ll=117) then grbp<="010";
	end if;
	if (ll=117 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=117 and cc>=98 and cc<100) then grbp<="010";
	end if;
	if (ll=117 and cc>=168 and cc<172) then grbp<="010";
	end if;
	if (cc=224 and ll=117) then grbp<="010";
	end if;
	if (ll=117 and cc>=224 and cc<227) then grbp<="010";
	end if;
	if (ll=117 and cc>=228 and cc<231) then grbp<="010";
	end if;
	if (cc=0 and ll=118) then grbp<="010";
	end if;
	if (ll=118 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=118 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=118 and cc>=63 and cc<89) then grbp<="010";
	end if;
	if (ll=118 and cc>=90 and cc<96) then grbp<="010";
	end if;
	if (ll=118 and cc>=97 and cc<100) then grbp<="010";
	end if;
	if (ll=118 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (ll=118 and cc>=223 and cc<231) then grbp<="010";
	end if;
	if (ll=119 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=119 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=119 and cc>=63 and cc<91) then grbp<="010";
	end if;
	if (ll=119 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=119 and cc>=97 and cc<99) then grbp<="010";
	end if;
	if (cc=223 and ll=119) then grbp<="010";
	end if;
	if (ll=119 and cc>=223 and cc<231) then grbp<="010";
	end if;
	if (ll=120 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=120 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=120 and cc>=63 and cc<90) then grbp<="010";
	end if;
	if (ll=120 and cc>=92 and cc<95) then grbp<="010";
	end if;
	if (ll=120 and cc>=96 and cc<100) then grbp<="010";
	end if;
	if (ll=120 and cc>=223 and cc<230) then grbp<="010";
	end if;
	if (ll=121 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=121 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=121 and cc>=63 and cc<87) then grbp<="010";
	end if;
	if (ll=121 and cc>=88 and cc<95) then grbp<="010";
	end if;
	if (ll=121 and cc>=96 and cc<101) then grbp<="010";
	end if;
	if (cc=223 and ll=121) then grbp<="010";
	end if;
	if (ll=121 and cc>=223 and cc<229) then grbp<="010";
	end if;
	if (ll=122 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=122 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=122 and cc>=63 and cc<87) then grbp<="010";
	end if;
	if (ll=122 and cc>=88 and cc<99) then grbp<="010";
	end if;
	if (cc=222 and ll=122) then grbp<="010";
	end if;
	if (ll=122 and cc>=222 and cc<224) then grbp<="010";
	end if;
	if (ll=122 and cc>=226 and cc<229) then grbp<="010";
	end if;
	if (ll=123 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=123 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=123 and cc>=63 and cc<93) then grbp<="010";
	end if;
	if (ll=123 and cc>=94 and cc<99) then grbp<="010";
	end if;
	if (ll=123 and cc>=103 and cc<105) then grbp<="010";
	end if;
	if (cc=222 and ll=123) then grbp<="010";
	end if;
	if (ll=123 and cc>=222 and cc<229) then grbp<="010";
	end if;
	if (ll=124 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=124 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=124 and cc>=63 and cc<88) then grbp<="010";
	end if;
	if (ll=124 and cc>=89 and cc<92) then grbp<="010";
	end if;
	if (ll=124 and cc>=93 and cc<100) then grbp<="010";
	end if;
	if (cc=104 and ll=124) then grbp<="010";
	end if;
	if (cc=113 and ll=124) then grbp<="010";
	end if;
	if (cc=203 and ll=124) then grbp<="010";
	end if;
	if (cc=221 and ll=124) then grbp<="010";
	end if;
	if (ll=124 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=124 and cc>=224 and cc<229) then grbp<="010";
	end if;
	if (ll=125 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=125 and cc>=27 and cc<59) then grbp<="010";
	end if;
	if (ll=125 and cc>=64 and cc<87) then grbp<="010";
	end if;
	if (ll=125 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=125 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=125 and cc>=97 and cc<100) then grbp<="010";
	end if;
	if (ll=125 and cc>=101 and cc<103) then grbp<="010";
	end if;
	if (cc=203 and ll=125) then grbp<="010";
	end if;
	if (cc=221 and ll=125) then grbp<="010";
	end if;
	if (ll=125 and cc>=221 and cc<228) then grbp<="010";
	end if;
	if (ll=126 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=126 and cc>=27 and cc<59) then grbp<="010";
	end if;
	if (ll=126 and cc>=63 and cc<91) then grbp<="010";
	end if;
	if (ll=126 and cc>=92 and cc<98) then grbp<="010";
	end if;
	if (ll=126 and cc>=101 and cc<104) then grbp<="010";
	end if;
	if (cc=221 and ll=126) then grbp<="010";
	end if;
	if (ll=126 and cc>=221 and cc<224) then grbp<="010";
	end if;
	if (ll=126 and cc>=225 and cc<228) then grbp<="010";
	end if;
	if (ll=127 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=127 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=127 and cc>=63 and cc<98) then grbp<="010";
	end if;
	if (ll=127 and cc>=100 and cc<104) then grbp<="010";
	end if;
	if (cc=221 and ll=127) then grbp<="010";
	end if;
	if (ll=127 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=127 and cc>=224 and cc<227) then grbp<="010";
	end if;
	if (ll=128 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=128 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=128 and cc>=64 and cc<90) then grbp<="010";
	end if;
	if (ll=128 and cc>=91 and cc<97) then grbp<="010";
	end if;
	if (ll=128 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (cc=221 and ll=128) then grbp<="010";
	end if;
	if (cc=224 and ll=128) then grbp<="010";
	end if;
	if (ll=128 and cc>=224 and cc<227) then grbp<="010";
	end if;
	if (ll=129 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=129 and cc>=27 and cc<59) then grbp<="010";
	end if;
	if (ll=129 and cc>=65 and cc<89) then grbp<="010";
	end if;
	if (ll=129 and cc>=90 and cc<97) then grbp<="010";
	end if;
	if (ll=129 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=129 and cc>=104 and cc<106) then grbp<="010";
	end if;
	if (cc=202 and ll=129) then grbp<="010";
	end if;
	if (cc=220 and ll=129) then grbp<="010";
	end if;
	if (ll=129 and cc>=220 and cc<223) then grbp<="010";
	end if;
	if (ll=129 and cc>=224 and cc<227) then grbp<="010";
	end if;
	if (ll=130 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=130 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (cc=65 and ll=130) then grbp<="010";
	end if;
	if (ll=130 and cc>=65 and cc<89) then grbp<="010";
	end if;
	if (ll=130 and cc>=90 and cc<101) then grbp<="010";
	end if;
	if (ll=130 and cc>=104 and cc<106) then grbp<="010";
	end if;
	if (cc=197 and ll=130) then grbp<="010";
	end if;
	if (cc=202 and ll=130) then grbp<="010";
	end if;
	if (cc=220 and ll=130) then grbp<="010";
	end if;
	if (ll=130 and cc>=220 and cc<226) then grbp<="010";
	end if;
	if (ll=131 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=131 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=131 and cc>=64 and cc<88) then grbp<="010";
	end if;
	if (ll=131 and cc>=89 and cc<95) then grbp<="010";
	end if;
	if (ll=131 and cc>=96 and cc<100) then grbp<="010";
	end if;
	if (ll=131 and cc>=102 and cc<106) then grbp<="010";
	end if;
	if (cc=132 and ll=131) then grbp<="010";
	end if;
	if (cc=196 and ll=131) then grbp<="010";
	end if;
	if (ll=131 and cc>=196 and cc<198) then grbp<="010";
	end if;
	if (ll=131 and cc>=219 and cc<226) then grbp<="010";
	end if;
	if (ll=132 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=132 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (cc=66 and ll=132) then grbp<="010";
	end if;
	if (ll=132 and cc>=66 and cc<95) then grbp<="010";
	end if;
	if (ll=132 and cc>=96 and cc<98) then grbp<="010";
	end if;
	if (cc=102 and ll=132) then grbp<="010";
	end if;
	if (cc=106 and ll=132) then grbp<="010";
	end if;
	if (ll=132 and cc>=106 and cc<108) then grbp<="010";
	end if;
	if (cc=218 and ll=132) then grbp<="010";
	end if;
	if (ll=132 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=132 and cc>=222 and cc<226) then grbp<="010";
	end if;
	if (ll=133 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=133 and cc>=27 and cc<58) then grbp<="010";
	end if;
	if (ll=133 and cc>=66 and cc<94) then grbp<="010";
	end if;
	if (ll=133 and cc>=95 and cc<99) then grbp<="010";
	end if;
	if (ll=133 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=133 and cc>=105 and cc<107) then grbp<="010";
	end if;
	if (cc=195 and ll=133) then grbp<="010";
	end if;
	if (ll=133 and cc>=195 and cc<197) then grbp<="010";
	end if;
	if (cc=218 and ll=133) then grbp<="010";
	end if;
	if (ll=133 and cc>=218 and cc<226) then grbp<="010";
	end if;
	if (ll=134 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=134 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=134 and cc>=65 and cc<99) then grbp<="010";
	end if;
	if (cc=105 and ll=134) then grbp<="010";
	end if;
	if (ll=134 and cc>=105 and cc<107) then grbp<="010";
	end if;
	if (cc=195 and ll=134) then grbp<="010";
	end if;
	if (ll=134 and cc>=195 and cc<197) then grbp<="010";
	end if;
	if (cc=218 and ll=134) then grbp<="010";
	end if;
	if (ll=134 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=134 and cc>=222 and cc<225) then grbp<="010";
	end if;
	if (ll=135 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=135 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=135 and cc>=64 and cc<102) then grbp<="010";
	end if;
	if (cc=107 and ll=135) then grbp<="010";
	end if;
	if (cc=111 and ll=135) then grbp<="010";
	end if;
	if (cc=126 and ll=135) then grbp<="010";
	end if;
	if (ll=135 and cc>=126 and cc<128) then grbp<="010";
	end if;
	if (ll=135 and cc>=194 and cc<196) then grbp<="010";
	end if;
	if (ll=135 and cc>=218 and cc<220) then grbp<="010";
	end if;
	if (ll=135 and cc>=221 and cc<225) then grbp<="010";
	end if;
	if (ll=136 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=136 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=66 and ll=136) then grbp<="010";
	end if;
	if (ll=136 and cc>=66 and cc<85) then grbp<="010";
	end if;
	if (ll=136 and cc>=86 and cc<102) then grbp<="010";
	end if;
	if (ll=136 and cc>=103 and cc<105) then grbp<="010";
	end if;
	if (cc=126 and ll=136) then grbp<="010";
	end if;
	if (cc=194 and ll=136) then grbp<="010";
	end if;
	if (cc=218 and ll=136) then grbp<="010";
	end if;
	if (ll=136 and cc>=218 and cc<220) then grbp<="010";
	end if;
	if (ll=136 and cc>=221 and cc<225) then grbp<="010";
	end if;
	if (ll=137 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=137 and cc>=27 and cc<58) then grbp<="010";
	end if;
	if (ll=137 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=137 and cc>=67 and cc<92) then grbp<="010";
	end if;
	if (ll=137 and cc>=93 and cc<100) then grbp<="010";
	end if;
	if (ll=137 and cc>=101 and cc<105) then grbp<="010";
	end if;
	if (ll=137 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (cc=115 and ll=137) then grbp<="010";
	end if;
	if (cc=124 and ll=137) then grbp<="010";
	end if;
	if (ll=137 and cc>=124 and cc<126) then grbp<="010";
	end if;
	if (cc=217 and ll=137) then grbp<="010";
	end if;
	if (ll=137 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=137 and cc>=221 and cc<224) then grbp<="010";
	end if;
	if (ll=138 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=138 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=67 and ll=138) then grbp<="010";
	end if;
	if (ll=138 and cc>=67 and cc<101) then grbp<="010";
	end if;
	if (ll=138 and cc>=102 and cc<105) then grbp<="010";
	end if;
	if (cc=113 and ll=138) then grbp<="010";
	end if;
	if (cc=192 and ll=138) then grbp<="010";
	end if;
	if (cc=196 and ll=138) then grbp<="010";
	end if;
	if (cc=200 and ll=138) then grbp<="010";
	end if;
	if (cc=217 and ll=138) then grbp<="010";
	end if;
	if (ll=138 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=138 and cc>=221 and cc<224) then grbp<="010";
	end if;
	if (ll=139 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=139 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=68 and ll=139) then grbp<="010";
	end if;
	if (ll=139 and cc>=68 and cc<101) then grbp<="010";
	end if;
	if (ll=139 and cc>=102 and cc<104) then grbp<="010";
	end if;
	if (cc=119 and ll=139) then grbp<="010";
	end if;
	if (cc=122 and ll=139) then grbp<="010";
	end if;
	if (cc=195 and ll=139) then grbp<="010";
	end if;
	if (ll=139 and cc>=195 and cc<197) then grbp<="010";
	end if;
	if (cc=217 and ll=139) then grbp<="010";
	end if;
	if (ll=139 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=139 and cc>=221 and cc<224) then grbp<="010";
	end if;
	if (ll=140 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=140 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=140 and cc>=67 and cc<104) then grbp<="010";
	end if;
	if (cc=118 and ll=140) then grbp<="010";
	end if;
	if (cc=120 and ll=140) then grbp<="010";
	end if;
	if (ll=140 and cc>=120 and cc<123) then grbp<="010";
	end if;
	if (cc=194 and ll=140) then grbp<="010";
	end if;
	if (ll=140 and cc>=194 and cc<197) then grbp<="010";
	end if;
	if (ll=140 and cc>=216 and cc<223) then grbp<="010";
	end if;
	if (ll=141 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=141 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=67 and ll=141) then grbp<="010";
	end if;
	if (ll=141 and cc>=67 and cc<98) then grbp<="010";
	end if;
	if (ll=141 and cc>=99 and cc<104) then grbp<="010";
	end if;
	if (ll=141 and cc>=120 and cc<123) then grbp<="010";
	end if;
	if (cc=190 and ll=141) then grbp<="010";
	end if;
	if (cc=192 and ll=141) then grbp<="010";
	end if;
	if (ll=141 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (ll=141 and cc>=216 and cc<218) then grbp<="010";
	end if;
	if (ll=141 and cc>=219 and cc<223) then grbp<="010";
	end if;
	if (ll=142 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=142 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=142 and cc>=67 and cc<99) then grbp<="010";
	end if;
	if (ll=142 and cc>=100 and cc<104) then grbp<="010";
	end if;
	if (ll=142 and cc>=107 and cc<114) then grbp<="010";
	end if;
	if (ll=142 and cc>=116 and cc<118) then grbp<="010";
	end if;
	if (ll=142 and cc>=119 and cc<123) then grbp<="010";
	end if;
	if (cc=140 and ll=142) then grbp<="010";
	end if;
	if (cc=146 and ll=142) then grbp<="010";
	end if;
	if (cc=191 and ll=142) then grbp<="010";
	end if;
	if (ll=142 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (ll=142 and cc>=216 and cc<218) then grbp<="010";
	end if;
	if (ll=142 and cc>=219 and cc<222) then grbp<="010";
	end if;
	if (ll=143 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=143 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=66 and ll=143) then grbp<="010";
	end if;
	if (cc=68 and ll=143) then grbp<="010";
	end if;
	if (ll=143 and cc>=68 and cc<102) then grbp<="010";
	end if;
	if (ll=143 and cc>=103 and cc<118) then grbp<="010";
	end if;
	if (cc=124 and ll=143) then grbp<="010";
	end if;
	if (cc=139 and ll=143) then grbp<="010";
	end if;
	if (ll=143 and cc>=139 and cc<141) then grbp<="010";
	end if;
	if (cc=146 and ll=143) then grbp<="010";
	end if;
	if (cc=190 and ll=143) then grbp<="010";
	end if;
	if (ll=143 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (cc=216 and ll=143) then grbp<="010";
	end if;
	if (ll=143 and cc>=216 and cc<222) then grbp<="010";
	end if;
	if (ll=144 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=144 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=144 and cc>=68 and cc<101) then grbp<="010";
	end if;
	if (ll=144 and cc>=103 and cc<108) then grbp<="010";
	end if;
	if (ll=144 and cc>=109 and cc<117) then grbp<="010";
	end if;
	if (ll=144 and cc>=123 and cc<126) then grbp<="010";
	end if;
	if (cc=189 and ll=144) then grbp<="010";
	end if;
	if (ll=144 and cc>=189 and cc<195) then grbp<="010";
	end if;
	if (cc=215 and ll=144) then grbp<="010";
	end if;
	if (ll=144 and cc>=215 and cc<222) then grbp<="010";
	end if;
	if (ll=145 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=145 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=67 and ll=145) then grbp<="010";
	end if;
	if (cc=69 and ll=145) then grbp<="010";
	end if;
	if (cc=71 and ll=145) then grbp<="010";
	end if;
	if (ll=145 and cc>=71 and cc<97) then grbp<="010";
	end if;
	if (ll=145 and cc>=98 and cc<103) then grbp<="010";
	end if;
	if (ll=145 and cc>=104 and cc<108) then grbp<="010";
	end if;
	if (ll=145 and cc>=109 and cc<117) then grbp<="010";
	end if;
	if (ll=145 and cc>=126 and cc<129) then grbp<="010";
	end if;
	if (cc=136 and ll=145) then grbp<="010";
	end if;
	if (cc=138 and ll=145) then grbp<="010";
	end if;
	if (cc=142 and ll=145) then grbp<="010";
	end if;
	if (cc=145 and ll=145) then grbp<="010";
	end if;
	if (cc=188 and ll=145) then grbp<="010";
	end if;
	if (ll=145 and cc>=188 and cc<195) then grbp<="010";
	end if;
	if (ll=145 and cc>=215 and cc<217) then grbp<="010";
	end if;
	if (cc=220 and ll=145) then grbp<="010";
	end if;
	if (ll=145 and cc>=220 and cc<222) then grbp<="010";
	end if;
	if (ll=146 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=146 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=146 and cc>=66 and cc<70) then grbp<="010";
	end if;
	if (ll=146 and cc>=71 and cc<101) then grbp<="010";
	end if;
	if (cc=105 and ll=146) then grbp<="010";
	end if;
	if (cc=109 and ll=146) then grbp<="010";
	end if;
	if (ll=146 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=146 and cc>=128 and cc<131) then grbp<="010";
	end if;
	if (cc=137 and ll=146) then grbp<="010";
	end if;
	if (cc=139 and ll=146) then grbp<="010";
	end if;
	if (ll=146 and cc>=139 and cc<141) then grbp<="010";
	end if;
	if (ll=146 and cc>=187 and cc<195) then grbp<="010";
	end if;
	if (cc=215 and ll=146) then grbp<="010";
	end if;
	if (ll=146 and cc>=215 and cc<222) then grbp<="010";
	end if;
	if (cc=0 and ll=147) then grbp<="010";
	end if;
	if (ll=147 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=147 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (cc=68 and ll=147) then grbp<="010";
	end if;
	if (cc=70 and ll=147) then grbp<="010";
	end if;
	if (cc=72 and ll=147) then grbp<="010";
	end if;
	if (ll=147 and cc>=72 and cc<102) then grbp<="010";
	end if;
	if (ll=147 and cc>=103 and cc<106) then grbp<="010";
	end if;
	if (ll=147 and cc>=107 and cc<116) then grbp<="010";
	end if;
	if (ll=147 and cc>=130 and cc<136) then grbp<="010";
	end if;
	if (ll=147 and cc>=186 and cc<194) then grbp<="010";
	end if;
	if (cc=218 and ll=147) then grbp<="010";
	end if;
	if (ll=147 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=148 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=148 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=148 and cc>=67 and cc<71) then grbp<="010";
	end if;
	if (ll=148 and cc>=72 and cc<102) then grbp<="010";
	end if;
	if (ll=148 and cc>=103 and cc<105) then grbp<="010";
	end if;
	if (ll=148 and cc>=107 and cc<113) then grbp<="010";
	end if;
	if (cc=185 and ll=148) then grbp<="010";
	end if;
	if (ll=148 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (ll=148 and cc>=214 and cc<217) then grbp<="010";
	end if;
	if (ll=148 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=149 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=149 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=149 and cc>=67 and cc<70) then grbp<="010";
	end if;
	if (ll=149 and cc>=71 and cc<115) then grbp<="010";
	end if;
	if (ll=149 and cc>=183 and cc<193) then grbp<="010";
	end if;
	if (cc=214 and ll=149) then grbp<="010";
	end if;
	if (ll=149 and cc>=214 and cc<221) then grbp<="010";
	end if;
	if (ll=150 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=150 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=150 and cc>=66 and cc<104) then grbp<="010";
	end if;
	if (ll=150 and cc>=105 and cc<114) then grbp<="010";
	end if;
	if (cc=122 and ll=150) then grbp<="010";
	end if;
	if (ll=150 and cc>=122 and cc<124) then grbp<="010";
	end if;
	if (ll=150 and cc>=181 and cc<192) then grbp<="010";
	end if;
	if (ll=150 and cc>=214 and cc<221) then grbp<="010";
	end if;
	if (ll=151 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=151 and cc>=28 and cc<58) then grbp<="010";
	end if;
	if (ll=151 and cc>=66 and cc<105) then grbp<="010";
	end if;
	if (ll=151 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=151 and cc>=110 and cc<112) then grbp<="010";
	end if;
	if (ll=151 and cc>=118 and cc<120) then grbp<="010";
	end if;
	if (cc=144 and ll=151) then grbp<="010";
	end if;
	if (cc=180 and ll=151) then grbp<="010";
	end if;
	if (ll=151 and cc>=180 and cc<191) then grbp<="010";
	end if;
	if (ll=151 and cc>=214 and cc<220) then grbp<="010";
	end if;
	if (ll=152 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=152 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=152 and cc>=67 and cc<106) then grbp<="010";
	end if;
	if (ll=152 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=121 and ll=152) then grbp<="010";
	end if;
	if (cc=126 and ll=152) then grbp<="010";
	end if;
	if (cc=179 and ll=152) then grbp<="010";
	end if;
	if (ll=152 and cc>=179 and cc<191) then grbp<="010";
	end if;
	if (ll=152 and cc>=213 and cc<219) then grbp<="010";
	end if;
	if (cc=0 and ll=153) then grbp<="010";
	end if;
	if (ll=153 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=153 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=153 and cc>=67 and cc<110) then grbp<="010";
	end if;
	if (ll=153 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (cc=142 and ll=153) then grbp<="010";
	end if;
	if (ll=153 and cc>=142 and cc<144) then grbp<="010";
	end if;
	if (ll=153 and cc>=177 and cc<190) then grbp<="010";
	end if;
	if (ll=153 and cc>=213 and cc<215) then grbp<="010";
	end if;
	if (ll=153 and cc>=216 and cc<219) then grbp<="010";
	end if;
	if (ll=154 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=154 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=154 and cc>=66 and cc<107) then grbp<="010";
	end if;
	if (cc=142 and ll=154) then grbp<="010";
	end if;
	if (cc=176 and ll=154) then grbp<="010";
	end if;
	if (ll=154 and cc>=176 and cc<189) then grbp<="010";
	end if;
	if (ll=154 and cc>=213 and cc<219) then grbp<="010";
	end if;
	if (ll=155 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=155 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=155 and cc>=66 and cc<70) then grbp<="010";
	end if;
	if (ll=155 and cc>=71 and cc<106) then grbp<="010";
	end if;
	if (cc=121 and ll=155) then grbp<="010";
	end if;
	if (cc=123 and ll=155) then grbp<="010";
	end if;
	if (cc=125 and ll=155) then grbp<="010";
	end if;
	if (cc=138 and ll=155) then grbp<="010";
	end if;
	if (cc=141 and ll=155) then grbp<="010";
	end if;
	if (ll=155 and cc>=141 and cc<143) then grbp<="010";
	end if;
	if (ll=155 and cc>=176 and cc<188) then grbp<="010";
	end if;
	if (cc=215 and ll=155) then grbp<="010";
	end if;
	if (ll=155 and cc>=215 and cc<218) then grbp<="010";
	end if;
	if (ll=156 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=156 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=156 and cc>=66 and cc<106) then grbp<="010";
	end if;
	if (cc=119 and ll=156) then grbp<="010";
	end if;
	if (cc=121 and ll=156) then grbp<="010";
	end if;
	if (ll=156 and cc>=121 and cc<123) then grbp<="010";
	end if;
	if (cc=140 and ll=156) then grbp<="010";
	end if;
	if (ll=156 and cc>=140 and cc<142) then grbp<="010";
	end if;
	if (ll=156 and cc>=175 and cc<187) then grbp<="010";
	end if;
	if (cc=212 and ll=156) then grbp<="010";
	end if;
	if (ll=156 and cc>=212 and cc<215) then grbp<="010";
	end if;
	if (ll=156 and cc>=216 and cc<218) then grbp<="010";
	end if;
	if (ll=157 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=157 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=157 and cc>=66 and cc<100) then grbp<="010";
	end if;
	if (ll=157 and cc>=101 and cc<107) then grbp<="010";
	end if;
	if (cc=120 and ll=157) then grbp<="010";
	end if;
	if (cc=124 and ll=157) then grbp<="010";
	end if;
	if (cc=126 and ll=157) then grbp<="010";
	end if;
	if (cc=139 and ll=157) then grbp<="010";
	end if;
	if (ll=157 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (cc=175 and ll=157) then grbp<="010";
	end if;
	if (ll=157 and cc>=175 and cc<186) then grbp<="010";
	end if;
	if (ll=157 and cc>=212 and cc<218) then grbp<="010";
	end if;
	if (ll=158 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=158 and cc>=28 and cc<59) then grbp<="010";
	end if;
	if (ll=158 and cc>=67 and cc<71) then grbp<="010";
	end if;
	if (ll=158 and cc>=72 and cc<100) then grbp<="010";
	end if;
	if (ll=158 and cc>=101 and cc<106) then grbp<="010";
	end if;
	if (cc=120 and ll=158) then grbp<="010";
	end if;
	if (cc=136 and ll=158) then grbp<="010";
	end if;
	if (cc=139 and ll=158) then grbp<="010";
	end if;
	if (ll=158 and cc>=139 and cc<141) then grbp<="010";
	end if;
	if (ll=158 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=158 and cc>=176 and cc<184) then grbp<="010";
	end if;
	if (ll=158 and cc>=212 and cc<218) then grbp<="010";
	end if;
	if (cc=0 and ll=159) then grbp<="010";
	end if;
	if (ll=159 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=159 and cc>=28 and cc<60) then grbp<="010";
	end if;
	if (ll=159 and cc>=67 and cc<72) then grbp<="010";
	end if;
	if (ll=159 and cc>=73 and cc<105) then grbp<="010";
	end if;
	if (cc=116 and ll=159) then grbp<="010";
	end if;
	if (cc=138 and ll=159) then grbp<="010";
	end if;
	if (ll=159 and cc>=138 and cc<140) then grbp<="010";
	end if;
	if (ll=159 and cc>=171 and cc<174) then grbp<="010";
	end if;
	if (ll=159 and cc>=176 and cc<182) then grbp<="010";
	end if;
	if (cc=211 and ll=159) then grbp<="010";
	end if;
	if (ll=159 and cc>=211 and cc<217) then grbp<="010";
	end if;
	if (ll=160 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=160 and cc>=28 and cc<60) then grbp<="010";
	end if;
	if (ll=160 and cc>=68 and cc<104) then grbp<="010";
	end if;
	if (cc=127 and ll=160) then grbp<="010";
	end if;
	if (cc=135 and ll=160) then grbp<="010";
	end if;
	if (cc=137 and ll=160) then grbp<="010";
	end if;
	if (ll=160 and cc>=137 and cc<139) then grbp<="010";
	end if;
	if (cc=172 and ll=160) then grbp<="010";
	end if;
	if (ll=160 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=160 and cc>=178 and cc<180) then grbp<="010";
	end if;
	if (ll=160 and cc>=211 and cc<217) then grbp<="010";
	end if;
	if (ll=161 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=161 and cc>=28 and cc<60) then grbp<="010";
	end if;
	if (ll=161 and cc>=69 and cc<92) then grbp<="010";
	end if;
	if (ll=161 and cc>=93 and cc<103) then grbp<="010";
	end if;
	if (ll=161 and cc>=117 and cc<119) then grbp<="010";
	end if;
	if (cc=134 and ll=161) then grbp<="010";
	end if;
	if (cc=137 and ll=161) then grbp<="010";
	end if;
	if (ll=161 and cc>=137 and cc<139) then grbp<="010";
	end if;
	if (ll=161 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (ll=161 and cc>=172 and cc<175) then grbp<="010";
	end if;
	if (cc=211 and ll=161) then grbp<="010";
	end if;
	if (ll=161 and cc>=211 and cc<215) then grbp<="010";
	end if;
	if (cc=0 and ll=162) then grbp<="010";
	end if;
	if (ll=162 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=162 and cc>=28 and cc<60) then grbp<="010";
	end if;
	if (ll=162 and cc>=69 and cc<102) then grbp<="010";
	end if;
	if (cc=117 and ll=162) then grbp<="010";
	end if;
	if (ll=162 and cc>=117 and cc<119) then grbp<="010";
	end if;
	if (cc=133 and ll=162) then grbp<="010";
	end if;
	if (cc=136 and ll=162) then grbp<="010";
	end if;
	if (ll=162 and cc>=136 and cc<138) then grbp<="010";
	end if;
	if (cc=170 and ll=162) then grbp<="010";
	end if;
	if (ll=162 and cc>=170 and cc<175) then grbp<="010";
	end if;
	if (ll=162 and cc>=211 and cc<217) then grbp<="010";
	end if;
	if (ll=163 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=163 and cc>=28 and cc<60) then grbp<="010";
	end if;
	if (cc=72 and ll=163) then grbp<="010";
	end if;
	if (ll=163 and cc>=72 and cc<101) then grbp<="010";
	end if;
	if (cc=124 and ll=163) then grbp<="010";
	end if;
	if (cc=135 and ll=163) then grbp<="010";
	end if;
	if (ll=163 and cc>=135 and cc<137) then grbp<="010";
	end if;
	if (ll=163 and cc>=170 and cc<175) then grbp<="010";
	end if;
	if (cc=211 and ll=163) then grbp<="010";
	end if;
	if (cc=213 and ll=163) then grbp<="010";
	end if;
	if (ll=163 and cc>=213 and cc<217) then grbp<="010";
	end if;
	if (ll=164 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=164 and cc>=28 and cc<61) then grbp<="010";
	end if;
	if (cc=72 and ll=164) then grbp<="010";
	end if;
	if (ll=164 and cc>=72 and cc<100) then grbp<="010";
	end if;
	if (cc=123 and ll=164) then grbp<="010";
	end if;
	if (cc=132 and ll=164) then grbp<="010";
	end if;
	if (cc=134 and ll=164) then grbp<="010";
	end if;
	if (ll=164 and cc>=134 and cc<137) then grbp<="010";
	end if;
	if (cc=170 and ll=164) then grbp<="010";
	end if;
	if (cc=172 and ll=164) then grbp<="010";
	end if;
	if (ll=164 and cc>=172 and cc<175) then grbp<="010";
	end if;
	if (cc=210 and ll=164) then grbp<="010";
	end if;
	if (ll=164 and cc>=210 and cc<216) then grbp<="010";
	end if;
	if (ll=165 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=165 and cc>=28 and cc<61) then grbp<="010";
	end if;
	if (ll=165 and cc>=70 and cc<100) then grbp<="010";
	end if;
	if (cc=133 and ll=165) then grbp<="010";
	end if;
	if (ll=165 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (cc=168 and ll=165) then grbp<="010";
	end if;
	if (ll=165 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (ll=165 and cc>=172 and cc<176) then grbp<="010";
	end if;
	if (ll=165 and cc>=210 and cc<216) then grbp<="010";
	end if;
	if (ll=166 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=166 and cc>=28 and cc<61) then grbp<="010";
	end if;
	if (ll=166 and cc>=71 and cc<98) then grbp<="010";
	end if;
	if (cc=121 and ll=166) then grbp<="010";
	end if;
	if (cc=133 and ll=166) then grbp<="010";
	end if;
	if (ll=166 and cc>=133 and cc<135) then grbp<="010";
	end if;
	if (cc=168 and ll=166) then grbp<="010";
	end if;
	if (ll=166 and cc>=168 and cc<170) then grbp<="010";
	end if;
	if (cc=175 and ll=166) then grbp<="010";
	end if;
	if (cc=178 and ll=166) then grbp<="010";
	end if;
	if (cc=187 and ll=166) then grbp<="010";
	end if;
	if (cc=210 and ll=166) then grbp<="010";
	end if;
	if (ll=166 and cc>=210 and cc<216) then grbp<="010";
	end if;
	if (ll=167 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=167 and cc>=28 and cc<61) then grbp<="010";
	end if;
	if (ll=167 and cc>=71 and cc<95) then grbp<="010";
	end if;
	if (cc=102 and ll=167) then grbp<="010";
	end if;
	if (cc=108 and ll=167) then grbp<="010";
	end if;
	if (ll=167 and cc>=108 and cc<110) then grbp<="010";
	end if;
	if (ll=167 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=167 and cc>=164 and cc<166) then grbp<="010";
	end if;
	if (ll=167 and cc>=168 and cc<172) then grbp<="010";
	end if;
	if (cc=175 and ll=167) then grbp<="010";
	end if;
	if (cc=178 and ll=167) then grbp<="010";
	end if;
	if (cc=186 and ll=167) then grbp<="010";
	end if;
	if (cc=209 and ll=167) then grbp<="010";
	end if;
	if (ll=167 and cc>=209 and cc<216) then grbp<="010";
	end if;
	if (ll=168 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=168 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (ll=168 and cc>=71 and cc<95) then grbp<="010";
	end if;
	if (ll=168 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (ll=168 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (ll=168 and cc>=164 and cc<168) then grbp<="010";
	end if;
	if (ll=168 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (ll=168 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=185 and ll=168) then grbp<="010";
	end if;
	if (cc=209 and ll=168) then grbp<="010";
	end if;
	if (ll=168 and cc>=209 and cc<215) then grbp<="010";
	end if;
	if (ll=169 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=169 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (ll=169 and cc>=71 and cc<98) then grbp<="010";
	end if;
	if (cc=114 and ll=169) then grbp<="010";
	end if;
	if (cc=131 and ll=169) then grbp<="010";
	end if;
	if (ll=169 and cc>=131 and cc<133) then grbp<="010";
	end if;
	if (ll=169 and cc>=164 and cc<173) then grbp<="010";
	end if;
	if (ll=169 and cc>=174 and cc<177) then grbp<="010";
	end if;
	if (ll=169 and cc>=209 and cc<215) then grbp<="010";
	end if;
	if (ll=170 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=170 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (ll=170 and cc>=71 and cc<88) then grbp<="010";
	end if;
	if (ll=170 and cc>=89 and cc<98) then grbp<="010";
	end if;
	if (cc=107 and ll=170) then grbp<="010";
	end if;
	if (cc=114 and ll=170) then grbp<="010";
	end if;
	if (ll=170 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (ll=170 and cc>=130 and cc<133) then grbp<="010";
	end if;
	if (ll=170 and cc>=164 and cc<169) then grbp<="010";
	end if;
	if (ll=170 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=170 and cc>=174 and cc<177) then grbp<="010";
	end if;
	if (cc=209 and ll=170) then grbp<="010";
	end if;
	if (ll=170 and cc>=209 and cc<215) then grbp<="010";
	end if;
	if (cc=0 and ll=171) then grbp<="010";
	end if;
	if (ll=171 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=171 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (ll=171 and cc>=70 and cc<83) then grbp<="010";
	end if;
	if (ll=171 and cc>=86 and cc<88) then grbp<="010";
	end if;
	if (ll=171 and cc>=89 and cc<98) then grbp<="010";
	end if;
	if (cc=107 and ll=171) then grbp<="010";
	end if;
	if (cc=114 and ll=171) then grbp<="010";
	end if;
	if (cc=131 and ll=171) then grbp<="010";
	end if;
	if (cc=165 and ll=171) then grbp<="010";
	end if;
	if (ll=171 and cc>=165 and cc<167) then grbp<="010";
	end if;
	if (ll=171 and cc>=168 and cc<173) then grbp<="010";
	end if;
	if (cc=183 and ll=171) then grbp<="010";
	end if;
	if (cc=208 and ll=171) then grbp<="010";
	end if;
	if (ll=171 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=172 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=172 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (ll=172 and cc>=70 and cc<83) then grbp<="010";
	end if;
	if (cc=91 and ll=172) then grbp<="010";
	end if;
	if (ll=172 and cc>=91 and cc<94) then grbp<="010";
	end if;
	if (ll=172 and cc>=95 and cc<98) then grbp<="010";
	end if;
	if (ll=172 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (cc=165 and ll=172) then grbp<="010";
	end if;
	if (ll=172 and cc>=165 and cc<169) then grbp<="010";
	end if;
	if (ll=172 and cc>=170 and cc<174) then grbp<="010";
	end if;
	if (cc=182 and ll=172) then grbp<="010";
	end if;
	if (cc=208 and ll=172) then grbp<="010";
	end if;
	if (ll=172 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=173 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=173 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=173 and cc>=70 and cc<86) then grbp<="010";
	end if;
	if (cc=92 and ll=173) then grbp<="010";
	end if;
	if (ll=173 and cc>=92 and cc<94) then grbp<="010";
	end if;
	if (cc=97 and ll=173) then grbp<="010";
	end if;
	if (ll=173 and cc>=97 and cc<101) then grbp<="010";
	end if;
	if (cc=118 and ll=173) then grbp<="010";
	end if;
	if (ll=173 and cc>=118 and cc<121) then grbp<="010";
	end if;
	if (cc=165 and ll=173) then grbp<="010";
	end if;
	if (ll=173 and cc>=165 and cc<170) then grbp<="010";
	end if;
	if (ll=173 and cc>=171 and cc<174) then grbp<="010";
	end if;
	if (cc=208 and ll=173) then grbp<="010";
	end if;
	if (ll=173 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=174 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=174 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=174 and cc>=70 and cc<87) then grbp<="010";
	end if;
	if (ll=174 and cc>=90 and cc<92) then grbp<="010";
	end if;
	if (ll=174 and cc>=96 and cc<101) then grbp<="010";
	end if;
	if (ll=174 and cc>=107 and cc<109) then grbp<="010";
	end if;
	if (ll=174 and cc>=165 and cc<169) then grbp<="010";
	end if;
	if (ll=174 and cc>=170 and cc<172) then grbp<="010";
	end if;
	if (ll=174 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=174 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=175 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=175 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=175 and cc>=70 and cc<92) then grbp<="010";
	end if;
	if (cc=99 and ll=175) then grbp<="010";
	end if;
	if (cc=108 and ll=175) then grbp<="010";
	end if;
	if (cc=166 and ll=175) then grbp<="010";
	end if;
	if (ll=175 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (cc=174 and ll=175) then grbp<="010";
	end if;
	if (cc=179 and ll=175) then grbp<="010";
	end if;
	if (ll=175 and cc>=179 and cc<182) then grbp<="010";
	end if;
	if (ll=175 and cc>=207 and cc<214) then grbp<="010";
	end if;
	if (ll=176 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=176 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=176 and cc>=71 and cc<92) then grbp<="010";
	end if;
	if (cc=108 and ll=176) then grbp<="010";
	end if;
	if (cc=166 and ll=176) then grbp<="010";
	end if;
	if (ll=176 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=176 and cc>=171 and cc<175) then grbp<="010";
	end if;
	if (ll=176 and cc>=179 and cc<182) then grbp<="010";
	end if;
	if (ll=176 and cc>=207 and cc<214) then grbp<="010";
	end if;
	if (ll=177 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=177 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=177 and cc>=71 and cc<92) then grbp<="010";
	end if;
	if (cc=110 and ll=177) then grbp<="010";
	end if;
	if (cc=124 and ll=177) then grbp<="010";
	end if;
	if (ll=177 and cc>=124 and cc<126) then grbp<="010";
	end if;
	if (ll=177 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=177 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=177 and cc>=179 and cc<182) then grbp<="010";
	end if;
	if (ll=177 and cc>=207 and cc<214) then grbp<="010";
	end if;
	if (ll=178 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=178 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=178 and cc>=70 and cc<93) then grbp<="010";
	end if;
	if (cc=123 and ll=178) then grbp<="010";
	end if;
	if (ll=178 and cc>=123 and cc<126) then grbp<="010";
	end if;
	if (ll=178 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=178 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=178 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=178 and cc>=207 and cc<213) then grbp<="010";
	end if;
	if (ll=179 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=179 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=179 and cc>=70 and cc<91) then grbp<="010";
	end if;
	if (cc=110 and ll=179) then grbp<="010";
	end if;
	if (cc=124 and ll=179) then grbp<="010";
	end if;
	if (ll=179 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=179 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (cc=175 and ll=179) then grbp<="010";
	end if;
	if (cc=179 and ll=179) then grbp<="010";
	end if;
	if (ll=179 and cc>=179 and cc<182) then grbp<="010";
	end if;
	if (ll=179 and cc>=207 and cc<213) then grbp<="010";
	end if;
	if (cc=0 and ll=180) then grbp<="010";
	end if;
	if (ll=180 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=180 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=180 and cc>=70 and cc<90) then grbp<="010";
	end if;
	if (cc=103 and ll=180) then grbp<="010";
	end if;
	if (cc=122 and ll=180) then grbp<="010";
	end if;
	if (ll=180 and cc>=122 and cc<126) then grbp<="010";
	end if;
	if (ll=180 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (cc=175 and ll=180) then grbp<="010";
	end if;
	if (cc=180 and ll=180) then grbp<="010";
	end if;
	if (cc=206 and ll=180) then grbp<="010";
	end if;
	if (ll=180 and cc>=206 and cc<213) then grbp<="010";
	end if;
	if (ll=181 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=181 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=181 and cc>=69 and cc<88) then grbp<="010";
	end if;
	if (cc=103 and ll=181) then grbp<="010";
	end if;
	if (cc=122 and ll=181) then grbp<="010";
	end if;
	if (ll=181 and cc>=122 and cc<126) then grbp<="010";
	end if;
	if (ll=181 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=181 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (cc=206 and ll=181) then grbp<="010";
	end if;
	if (ll=181 and cc>=206 and cc<212) then grbp<="010";
	end if;
	if (ll=182 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=182 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=182 and cc>=69 and cc<88) then grbp<="010";
	end if;
	if (cc=103 and ll=182) then grbp<="010";
	end if;
	if (cc=121 and ll=182) then grbp<="010";
	end if;
	if (ll=182 and cc>=121 and cc<125) then grbp<="010";
	end if;
	if (ll=182 and cc>=167 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=182) then grbp<="010";
	end if;
	if (cc=206 and ll=182) then grbp<="010";
	end if;
	if (ll=182 and cc>=206 and cc<212) then grbp<="010";
	end if;
	if (cc=250 and ll=182) then grbp<="010";
	end if;
	if (cc=0 and ll=183) then grbp<="010";
	end if;
	if (ll=183 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=183 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=183 and cc>=69 and cc<88) then grbp<="010";
	end if;
	if (ll=183 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=183 and cc>=122 and cc<125) then grbp<="010";
	end if;
	if (ll=183 and cc>=167 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=183) then grbp<="010";
	end if;
	if (cc=205 and ll=183) then grbp<="010";
	end if;
	if (ll=183 and cc>=205 and cc<212) then grbp<="010";
	end if;
	if (cc=250 and ll=183) then grbp<="010";
	end if;
	if (cc=0 and ll=184) then grbp<="010";
	end if;
	if (ll=184 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=184 and cc>=28 and cc<64) then grbp<="010";
	end if;
	if (ll=184 and cc>=68 and cc<88) then grbp<="010";
	end if;
	if (cc=120 and ll=184) then grbp<="010";
	end if;
	if (cc=122 and ll=184) then grbp<="010";
	end if;
	if (ll=184 and cc>=122 and cc<124) then grbp<="010";
	end if;
	if (ll=184 and cc>=167 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=184) then grbp<="010";
	end if;
	if (cc=205 and ll=184) then grbp<="010";
	end if;
	if (ll=184 and cc>=205 and cc<211) then grbp<="010";
	end if;
	if (cc=0 and ll=185) then grbp<="010";
	end if;
	if (ll=185 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=185 and cc>=29 and cc<65) then grbp<="010";
	end if;
	if (ll=185 and cc>=68 and cc<88) then grbp<="010";
	end if;
	if (cc=119 and ll=185) then grbp<="010";
	end if;
	if (cc=121 and ll=185) then grbp<="010";
	end if;
	if (ll=185 and cc>=121 and cc<123) then grbp<="010";
	end if;
	if (ll=185 and cc>=167 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=185) then grbp<="010";
	end if;
	if (cc=205 and ll=185) then grbp<="010";
	end if;
	if (ll=185 and cc>=205 and cc<211) then grbp<="010";
	end if;
	if (cc=0 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=186 and cc>=28 and cc<65) then grbp<="010";
	end if;
	if (ll=186 and cc>=68 and cc<85) then grbp<="010";
	end if;
	if (ll=186 and cc>=90 and cc<92) then grbp<="010";
	end if;
	if (cc=121 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=121 and cc<123) then grbp<="010";
	end if;
	if (cc=167 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=186) then grbp<="010";
	end if;
	if (cc=205 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=205 and cc<211) then grbp<="010";
	end if;
	if (cc=0 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=187 and cc>=28 and cc<55) then grbp<="010";
	end if;
	if (ll=187 and cc>=56 and cc<65) then grbp<="010";
	end if;
	if (ll=187 and cc>=68 and cc<82) then grbp<="010";
	end if;
	if (cc=86 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=86 and cc<88) then grbp<="010";
	end if;
	if (cc=106 and ll=187) then grbp<="010";
	end if;
	if (cc=118 and ll=187) then grbp<="010";
	end if;
	if (cc=120 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=120 and cc<122) then grbp<="010";
	end if;
	if (cc=167 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=205 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=205 and cc<210) then grbp<="010";
	end if;
	if (cc=0 and ll=188) then grbp<="010";
	end if;
	if (ll=188 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=188 and cc>=28 and cc<54) then grbp<="010";
	end if;
	if (ll=188 and cc>=55 and cc<65) then grbp<="010";
	end if;
	if (ll=188 and cc>=68 and cc<83) then grbp<="010";
	end if;
	if (cc=106 and ll=188) then grbp<="010";
	end if;
	if (ll=188 and cc>=106 and cc<108) then grbp<="010";
	end if;
	if (ll=188 and cc>=118 and cc<122) then grbp<="010";
	end if;
	if (cc=168 and ll=188) then grbp<="010";
	end if;
	if (ll=188 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=205 and ll=188) then grbp<="010";
	end if;
	if (ll=188 and cc>=205 and cc<210) then grbp<="010";
	end if;
	if (cc=222 and ll=188) then grbp<="010";
	end if;
	if (cc=250 and ll=188) then grbp<="010";
	end if;
	if (cc=0 and ll=189) then grbp<="010";
	end if;
	if (ll=189 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=189 and cc>=28 and cc<54) then grbp<="010";
	end if;
	if (ll=189 and cc>=55 and cc<66) then grbp<="010";
	end if;
	if (ll=189 and cc>=68 and cc<85) then grbp<="010";
	end if;
	if (cc=117 and ll=189) then grbp<="010";
	end if;
	if (cc=119 and ll=189) then grbp<="010";
	end if;
	if (ll=189 and cc>=119 and cc<121) then grbp<="010";
	end if;
	if (ll=189 and cc>=141 and cc<143) then grbp<="010";
	end if;
	if (ll=189 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=204 and ll=189) then grbp<="010";
	end if;
	if (ll=189 and cc>=204 and cc<210) then grbp<="010";
	end if;
	if (cc=250 and ll=189) then grbp<="010";
	end if;
	if (cc=0 and ll=190) then grbp<="010";
	end if;
	if (ll=190 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=190 and cc>=28 and cc<66) then grbp<="010";
	end if;
	if (ll=190 and cc>=68 and cc<84) then grbp<="010";
	end if;
	if (cc=107 and ll=190) then grbp<="010";
	end if;
	if (cc=117 and ll=190) then grbp<="010";
	end if;
	if (ll=190 and cc>=117 and cc<121) then grbp<="010";
	end if;
	if (cc=168 and ll=190) then grbp<="010";
	end if;
	if (ll=190 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=204 and ll=190) then grbp<="010";
	end if;
	if (ll=190 and cc>=204 and cc<210) then grbp<="010";
	end if;
	if (cc=250 and ll=190) then grbp<="010";
	end if;
	if (cc=0 and ll=191) then grbp<="010";
	end if;
	if (ll=191 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=191 and cc>=28 and cc<66) then grbp<="010";
	end if;
	if (ll=191 and cc>=68 and cc<83) then grbp<="010";
	end if;
	if (cc=107 and ll=191) then grbp<="010";
	end if;
	if (ll=191 and cc>=107 and cc<109) then grbp<="010";
	end if;
	if (cc=118 and ll=191) then grbp<="010";
	end if;
	if (ll=191 and cc>=118 and cc<120) then grbp<="010";
	end if;
	if (cc=168 and ll=191) then grbp<="010";
	end if;
	if (ll=191 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (ll=191 and cc>=176 and cc<178) then grbp<="010";
	end if;
	if (cc=204 and ll=191) then grbp<="010";
	end if;
	if (ll=191 and cc>=204 and cc<209) then grbp<="010";
	end if;
	if (cc=223 and ll=191) then grbp<="010";
	end if;
	if (cc=228 and ll=191) then grbp<="010";
	end if;
	if (cc=248 and ll=191) then grbp<="010";
	end if;
	if (cc=250 and ll=191) then grbp<="010";
	end if;
	if (cc=0 and ll=192) then grbp<="010";
	end if;
	if (ll=192 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=192 and cc>=28 and cc<66) then grbp<="010";
	end if;
	if (ll=192 and cc>=68 and cc<83) then grbp<="010";
	end if;
	if (cc=111 and ll=192) then grbp<="010";
	end if;
	if (cc=116 and ll=192) then grbp<="010";
	end if;
	if (ll=192 and cc>=116 and cc<120) then grbp<="010";
	end if;
	if (cc=168 and ll=192) then grbp<="010";
	end if;
	if (ll=192 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (ll=192 and cc>=176 and cc<178) then grbp<="010";
	end if;
	if (ll=192 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=192 and cc>=203 and cc<209) then grbp<="010";
	end if;
	if (cc=227 and ll=192) then grbp<="010";
	end if;
	if (ll=192 and cc>=227 and cc<229) then grbp<="010";
	end if;
	if (cc=250 and ll=192) then grbp<="010";
	end if;
	if (cc=0 and ll=193) then grbp<="010";
	end if;
	if (ll=193 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=193 and cc>=28 and cc<67) then grbp<="010";
	end if;
	if (ll=193 and cc>=69 and cc<82) then grbp<="010";
	end if;
	if (cc=115 and ll=193) then grbp<="010";
	end if;
	if (cc=117 and ll=193) then grbp<="010";
	end if;
	if (ll=193 and cc>=117 and cc<119) then grbp<="010";
	end if;
	if (ll=193 and cc>=138 and cc<140) then grbp<="010";
	end if;
	if (ll=193 and cc>=168 and cc<172) then grbp<="010";
	end if;
	if (cc=180 and ll=193) then grbp<="010";
	end if;
	if (ll=193 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=193 and cc>=203 and cc<209) then grbp<="010";
	end if;
	if (cc=228 and ll=193) then grbp<="010";
	end if;
	if (ll=193 and cc>=228 and cc<233) then grbp<="010";
	end if;
	if (cc=0 and ll=194) then grbp<="010";
	end if;
	if (ll=194 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=194 and cc>=28 and cc<67) then grbp<="010";
	end if;
	if (ll=194 and cc>=69 and cc<81) then grbp<="010";
	end if;
	if (ll=194 and cc>=115 and cc<119) then grbp<="010";
	end if;
	if (cc=168 and ll=194) then grbp<="010";
	end if;
	if (ll=194 and cc>=168 and cc<172) then grbp<="010";
	end if;
	if (ll=194 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=194 and cc>=203 and cc<209) then grbp<="010";
	end if;
	if (cc=230 and ll=194) then grbp<="010";
	end if;
	if (cc=232 and ll=194) then grbp<="010";
	end if;
	if (cc=234 and ll=194) then grbp<="010";
	end if;
	if (cc=250 and ll=194) then grbp<="010";
	end if;
	if (cc=0 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=195 and cc>=28 and cc<67) then grbp<="010";
	end if;
	if (ll=195 and cc>=68 and cc<80) then grbp<="010";
	end if;
	if (cc=116 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=116 and cc<118) then grbp<="010";
	end if;
	if (cc=168 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=168 and cc<172) then grbp<="010";
	end if;
	if (cc=203 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=203 and cc<209) then grbp<="010";
	end if;
	if (cc=232 and ll=195) then grbp<="010";
	end if;
	if (cc=234 and ll=195) then grbp<="010";
	end if;
	if (cc=236 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=236 and cc<238) then grbp<="010";
	end if;
	if (cc=244 and ll=195) then grbp<="010";
	end if;
	if (cc=249 and ll=195) then grbp<="010";
	end if;
	if (ll=195 and cc>=249 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=196) then grbp<="010";
	end if;
	if (ll=196 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=196 and cc>=29 and cc<75) then grbp<="010";
	end if;
	if (ll=196 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (cc=114 and ll=196) then grbp<="010";
	end if;
	if (cc=116 and ll=196) then grbp<="010";
	end if;
	if (ll=196 and cc>=116 and cc<118) then grbp<="010";
	end if;
	if (ll=196 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=180 and ll=196) then grbp<="010";
	end if;
	if (cc=202 and ll=196) then grbp<="010";
	end if;
	if (ll=196 and cc>=202 and cc<209) then grbp<="010";
	end if;
	if (ll=196 and cc>=229 and cc<231) then grbp<="010";
	end if;
	if (ll=196 and cc>=234 and cc<237) then grbp<="010";
	end if;
	if (ll=196 and cc>=238 and cc<241) then grbp<="010";
	end if;
	if (cc=0 and ll=197) then grbp<="010";
	end if;
	if (ll=197 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=197 and cc>=29 and cc<74) then grbp<="010";
	end if;
	if (ll=197 and cc>=77 and cc<79) then grbp<="010";
	end if;
	if (cc=113 and ll=197) then grbp<="010";
	end if;
	if (ll=197 and cc>=113 and cc<117) then grbp<="010";
	end if;
	if (ll=197 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (ll=197 and cc>=177 and cc<179) then grbp<="010";
	end if;
	if (ll=197 and cc>=180 and cc<182) then grbp<="010";
	end if;
	if (ll=197 and cc>=202 and cc<208) then grbp<="010";
	end if;
	if (cc=233 and ll=197) then grbp<="010";
	end if;
	if (ll=197 and cc>=233 and cc<236) then grbp<="010";
	end if;
	if (ll=197 and cc>=237 and cc<242) then grbp<="010";
	end if;
	if (cc=0 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=198 and cc>=28 and cc<73) then grbp<="010";
	end if;
	if (ll=198 and cc>=77 and cc<79) then grbp<="010";
	end if;
	if (cc=101 and ll=198) then grbp<="010";
	end if;
	if (cc=113 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=113 and cc<117) then grbp<="010";
	end if;
	if (cc=169 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (ll=198 and cc>=177 and cc<179) then grbp<="010";
	end if;
	if (cc=202 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=202 and cc<208) then grbp<="010";
	end if;
	if (cc=237 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=237 and cc<244) then grbp<="010";
	end if;
	if (ll=199 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=199 and cc>=28 and cc<72) then grbp<="010";
	end if;
	if (ll=199 and cc>=75 and cc<79) then grbp<="010";
	end if;
	if (cc=104 and ll=199) then grbp<="010";
	end if;
	if (cc=114 and ll=199) then grbp<="010";
	end if;
	if (ll=199 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (cc=169 and ll=199) then grbp<="010";
	end if;
	if (ll=199 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (ll=199 and cc>=177 and cc<179) then grbp<="010";
	end if;
	if (cc=202 and ll=199) then grbp<="010";
	end if;
	if (ll=199 and cc>=202 and cc<208) then grbp<="010";
	end if;
	if (ll=199 and cc>=234 and cc<240) then grbp<="010";
	end if;
	if (ll=199 and cc>=241 and cc<244) then grbp<="010";
	end if;
	if (ll=200 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=200 and cc>=28 and cc<68) then grbp<="010";
	end if;
	if (ll=200 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (ll=200 and cc>=74 and cc<79) then grbp<="010";
	end if;
	if (cc=112 and ll=200) then grbp<="010";
	end if;
	if (ll=200 and cc>=112 and cc<116) then grbp<="010";
	end if;
	if (ll=200 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (ll=200 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=200) then grbp<="010";
	end if;
	if (cc=202 and ll=200) then grbp<="010";
	end if;
	if (ll=200 and cc>=202 and cc<208) then grbp<="010";
	end if;
	if (ll=200 and cc>=232 and cc<234) then grbp<="010";
	end if;
	if (ll=200 and cc>=235 and cc<239) then grbp<="010";
	end if;
	if (ll=200 and cc>=240 and cc<249) then grbp<="010";
	end if;
	if (ll=201 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=201 and cc>=28 and cc<65) then grbp<="010";
	end if;
	if (ll=201 and cc>=66 and cc<68) then grbp<="010";
	end if;
	if (cc=74 and ll=201) then grbp<="010";
	end if;
	if (ll=201 and cc>=74 and cc<78) then grbp<="010";
	end if;
	if (cc=91 and ll=201) then grbp<="010";
	end if;
	if (ll=201 and cc>=91 and cc<93) then grbp<="010";
	end if;
	if (ll=201 and cc>=113 and cc<115) then grbp<="010";
	end if;
	if (ll=201 and cc>=131 and cc<135) then grbp<="010";
	end if;
	if (ll=201 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (cc=181 and ll=201) then grbp<="010";
	end if;
	if (cc=201 and ll=201) then grbp<="010";
	end if;
	if (ll=201 and cc>=201 and cc<207) then grbp<="010";
	end if;
	if (ll=201 and cc>=234 and cc<245) then grbp<="010";
	end if;
	if (ll=201 and cc>=246 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=202 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (ll=202 and cc>=64 and cc<71) then grbp<="010";
	end if;
	if (ll=202 and cc>=73 and cc<78) then grbp<="010";
	end if;
	if (cc=113 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=113 and cc<115) then grbp<="010";
	end if;
	if (ll=202 and cc>=130 and cc<137) then grbp<="010";
	end if;
	if (ll=202 and cc>=169 and cc<172) then grbp<="010";
	end if;
	if (ll=202 and cc>=177 and cc<179) then grbp<="010";
	end if;
	if (cc=201 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=201 and cc<207) then grbp<="010";
	end if;
	if (cc=237 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=237 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=203) then grbp<="010";
	end if;
	if (ll=203 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=203 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (cc=69 and ll=203) then grbp<="010";
	end if;
	if (cc=72 and ll=203) then grbp<="010";
	end if;
	if (ll=203 and cc>=72 and cc<77) then grbp<="010";
	end if;
	if (ll=203 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=203 and cc>=129 and cc<138) then grbp<="010";
	end if;
	if (ll=203 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (cc=181 and ll=203) then grbp<="010";
	end if;
	if (cc=201 and ll=203) then grbp<="010";
	end if;
	if (ll=203 and cc>=201 and cc<207) then grbp<="010";
	end if;
	if (ll=203 and cc>=241 and cc<244) then grbp<="010";
	end if;
	if (ll=203 and cc>=245 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=204 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (ll=204 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (cc=72 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=72 and cc<77) then grbp<="010";
	end if;
	if (cc=104 and ll=204) then grbp<="010";
	end if;
	if (cc=110 and ll=204) then grbp<="010";
	end if;
	if (cc=112 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=204 and cc>=128 and cc<140) then grbp<="010";
	end if;
	if (ll=204 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=181 and ll=204) then grbp<="010";
	end if;
	if (cc=201 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=201 and cc<207) then grbp<="010";
	end if;
	if (cc=240 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=240 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=205) then grbp<="010";
	end if;
	if (ll=205 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=205 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (cc=69 and ll=205) then grbp<="010";
	end if;
	if (cc=73 and ll=205) then grbp<="010";
	end if;
	if (ll=205 and cc>=73 and cc<76) then grbp<="010";
	end if;
	if (ll=205 and cc>=110 and cc<114) then grbp<="010";
	end if;
	if (ll=205 and cc>=128 and cc<141) then grbp<="010";
	end if;
	if (ll=205 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=201 and ll=205) then grbp<="010";
	end if;
	if (ll=205 and cc>=201 and cc<206) then grbp<="010";
	end if;
	if (ll=205 and cc>=241 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=206 and cc>=29 and cc<62) then grbp<="010";
	end if;
	if (cc=73 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=73 and cc<76) then grbp<="010";
	end if;
	if (cc=101 and ll=206) then grbp<="010";
	end if;
	if (cc=111 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=206 and cc>=127 and cc<142) then grbp<="010";
	end if;
	if (ll=206 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=200 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=200 and cc<206) then grbp<="010";
	end if;
	if (ll=206 and cc>=241 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=207 and cc>=28 and cc<62) then grbp<="010";
	end if;
	if (cc=71 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (cc=83 and ll=207) then grbp<="010";
	end if;
	if (cc=109 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=109 and cc<112) then grbp<="010";
	end if;
	if (ll=207 and cc>=126 and cc<143) then grbp<="010";
	end if;
	if (ll=207 and cc>=164 and cc<172) then grbp<="010";
	end if;
	if (cc=200 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=200 and cc<206) then grbp<="010";
	end if;
	if (ll=207 and cc>=242 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=208) then grbp<="010";
	end if;
	if (ll=208 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=208 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (cc=70 and ll=208) then grbp<="010";
	end if;
	if (ll=208 and cc>=70 and cc<74) then grbp<="010";
	end if;
	if (cc=109 and ll=208) then grbp<="010";
	end if;
	if (ll=208 and cc>=109 and cc<112) then grbp<="010";
	end if;
	if (ll=208 and cc>=126 and cc<132) then grbp<="010";
	end if;
	if (ll=208 and cc>=134 and cc<144) then grbp<="010";
	end if;
	if (ll=208 and cc>=163 and cc<173) then grbp<="010";
	end if;
	if (ll=208 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=208 and cc>=200 and cc<206) then grbp<="010";
	end if;
	if (ll=208 and cc>=244 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=209) then grbp<="010";
	end if;
	if (ll=209 and cc>=0 and cc<18) then grbp<="010";
	end if;
	if (ll=209 and cc>=28 and cc<63) then grbp<="010";
	end if;
	if (ll=209 and cc>=70 and cc<75) then grbp<="010";
	end if;
	if (cc=108 and ll=209) then grbp<="010";
	end if;
	if (cc=110 and ll=209) then grbp<="010";
	end if;
	if (ll=209 and cc>=110 and cc<112) then grbp<="010";
	end if;
	if (ll=209 and cc>=125 and cc<133) then grbp<="010";
	end if;
	if (ll=209 and cc>=134 and cc<145) then grbp<="010";
	end if;
	if (ll=209 and cc>=162 and cc<173) then grbp<="010";
	end if;
	if (ll=209 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=209 and cc>=200 and cc<206) then grbp<="010";
	end if;
	if (ll=209 and cc>=244 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=210 and cc>=29 and cc<59) then grbp<="010";
	end if;
	if (ll=210 and cc>=60 and cc<63) then grbp<="010";
	end if;
	if (cc=66 and ll=210) then grbp<="010";
	end if;
	if (cc=70 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=70 and cc<74) then grbp<="010";
	end if;
	if (cc=94 and ll=210) then grbp<="010";
	end if;
	if (cc=103 and ll=210) then grbp<="010";
	end if;
	if (cc=108 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (ll=210 and cc>=124 and cc<134) then grbp<="010";
	end if;
	if (ll=210 and cc>=135 and cc<145) then grbp<="010";
	end if;
	if (ll=210 and cc>=161 and cc<173) then grbp<="010";
	end if;
	if (cc=181 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=210 and cc>=200 and cc<205) then grbp<="010";
	end if;
	if (ll=210 and cc>=245 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=211 and cc>=29 and cc<59) then grbp<="010";
	end if;
	if (ll=211 and cc>=60 and cc<63) then grbp<="010";
	end if;
	if (cc=67 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (cc=94 and ll=211) then grbp<="010";
	end if;
	if (cc=109 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=109 and cc<111) then grbp<="010";
	end if;
	if (ll=211 and cc>=123 and cc<146) then grbp<="010";
	end if;
	if (cc=160 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=160 and cc<173) then grbp<="010";
	end if;
	if (cc=181 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=211 and cc>=199 and cc<205) then grbp<="010";
	end if;
	if (ll=211 and cc>=246 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=212 and cc>=29 and cc<59) then grbp<="010";
	end if;
	if (ll=212 and cc>=61 and cc<63) then grbp<="010";
	end if;
	if (ll=212 and cc>=67 and cc<72) then grbp<="010";
	end if;
	if (cc=86 and ll=212) then grbp<="010";
	end if;
	if (cc=94 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=94 and cc<96) then grbp<="010";
	end if;
	if (cc=109 and ll=212) then grbp<="010";
	end if;
	if (cc=123 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=123 and cc<132) then grbp<="010";
	end if;
	if (ll=212 and cc>=133 and cc<135) then grbp<="010";
	end if;
	if (ll=212 and cc>=136 and cc<148) then grbp<="010";
	end if;
	if (ll=212 and cc>=160 and cc<174) then grbp<="010";
	end if;
	if (cc=181 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=212 and cc>=199 and cc<205) then grbp<="010";
	end if;
	if (cc=247 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=247 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=213 and cc>=29 and cc<56) then grbp<="010";
	end if;
	if (ll=213 and cc>=57 and cc<59) then grbp<="010";
	end if;
	if (cc=65 and ll=213) then grbp<="010";
	end if;
	if (cc=67 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=67 and cc<69) then grbp<="010";
	end if;
	if (cc=107 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=107 and cc<110) then grbp<="010";
	end if;
	if (ll=213 and cc>=122 and cc<130) then grbp<="010";
	end if;
	if (cc=137 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=137 and cc<148) then grbp<="010";
	end if;
	if (cc=160 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=160 and cc<164) then grbp<="010";
	end if;
	if (ll=213 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (cc=181 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (ll=213 and cc>=199 and cc<205) then grbp<="010";
	end if;
	if (cc=245 and ll=213) then grbp<="010";
	end if;
	if (cc=247 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=247 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=0 and cc<18) then grbp<="010";
	end if;
	if (ll=214 and cc>=29 and cc<54) then grbp<="010";
	end if;
	if (ll=214 and cc>=57 and cc<69) then grbp<="010";
	end if;
	if (cc=80 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=80 and cc<82) then grbp<="010";
	end if;
	if (ll=214 and cc>=108 and cc<110) then grbp<="010";
	end if;
	if (ll=214 and cc>=121 and cc<126) then grbp<="010";
	end if;
	if (ll=214 and cc>=138 and cc<149) then grbp<="010";
	end if;
	if (ll=214 and cc>=159 and cc<162) then grbp<="010";
	end if;
	if (ll=214 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (cc=181 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=181 and cc<184) then grbp<="010";
	end if;
	if (ll=214 and cc>=199 and cc<205) then grbp<="010";
	end if;
	if (cc=243 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=243 and cc<245) then grbp<="010";
	end if;
	if (ll=214 and cc>=246 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=215) then grbp<="010";
	end if;
	if (ll=215 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=215 and cc>=29 and cc<54) then grbp<="010";
	end if;
	if (ll=215 and cc>=56 and cc<62) then grbp<="010";
	end if;
	if (ll=215 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (cc=77 and ll=215) then grbp<="010";
	end if;
	if (cc=85 and ll=215) then grbp<="010";
	end if;
	if (cc=95 and ll=215) then grbp<="010";
	end if;
	if (cc=106 and ll=215) then grbp<="010";
	end if;
	if (cc=108 and ll=215) then grbp<="010";
	end if;
	if (cc=121 and ll=215) then grbp<="010";
	end if;
	if (ll=215 and cc>=121 and cc<125) then grbp<="010";
	end if;
	if (ll=215 and cc>=139 and cc<149) then grbp<="010";
	end if;
	if (cc=179 and ll=215) then grbp<="010";
	end if;
	if (cc=181 and ll=215) then grbp<="010";
	end if;
	if (ll=215 and cc>=181 and cc<184) then grbp<="010";
	end if;
	if (ll=215 and cc>=199 and cc<205) then grbp<="010";
	end if;
	if (ll=215 and cc>=242 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=216 and cc>=28 and cc<53) then grbp<="010";
	end if;
	if (ll=216 and cc>=56 and cc<66) then grbp<="010";
	end if;
	if (cc=76 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=76 and cc<78) then grbp<="010";
	end if;
	if (cc=106 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=216 and cc>=120 and cc<123) then grbp<="010";
	end if;
	if (cc=140 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=140 and cc<149) then grbp<="010";
	end if;
	if (ll=216 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (cc=182 and ll=216) then grbp<="010";
	end if;
	if (cc=199 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=199 and cc<204) then grbp<="010";
	end if;
	if (cc=242 and ll=216) then grbp<="010";
	end if;
	if (cc=244 and ll=216) then grbp<="010";
	end if;
	if (ll=216 and cc>=244 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=217 and cc>=28 and cc<53) then grbp<="010";
	end if;
	if (ll=217 and cc>=56 and cc<61) then grbp<="010";
	end if;
	if (ll=217 and cc>=62 and cc<65) then grbp<="010";
	end if;
	if (cc=107 and ll=217) then grbp<="010";
	end if;
	if (cc=120 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=120 and cc<123) then grbp<="010";
	end if;
	if (cc=135 and ll=217) then grbp<="010";
	end if;
	if (cc=140 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=217 and cc>=157 and cc<159) then grbp<="010";
	end if;
	if (ll=217 and cc>=164 and cc<166) then grbp<="010";
	end if;
	if (cc=182 and ll=217) then grbp<="010";
	end if;
	if (cc=199 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=199 and cc<204) then grbp<="010";
	end if;
	if (ll=217 and cc>=240 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=218) then grbp<="010";
	end if;
	if (ll=218 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=218 and cc>=28 and cc<52) then grbp<="010";
	end if;
	if (ll=218 and cc>=56 and cc<60) then grbp<="010";
	end if;
	if (ll=218 and cc>=61 and cc<65) then grbp<="010";
	end if;
	if (cc=105 and ll=218) then grbp<="010";
	end if;
	if (ll=218 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=218 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (cc=136 and ll=218) then grbp<="010";
	end if;
	if (cc=141 and ll=218) then grbp<="010";
	end if;
	if (ll=218 and cc>=141 and cc<150) then grbp<="010";
	end if;
	if (cc=163 and ll=218) then grbp<="010";
	end if;
	if (cc=165 and ll=218) then grbp<="010";
	end if;
	if (ll=218 and cc>=165 and cc<167) then grbp<="010";
	end if;
	if (cc=182 and ll=218) then grbp<="010";
	end if;
	if (ll=218 and cc>=182 and cc<184) then grbp<="010";
	end if;
	if (ll=218 and cc>=198 and cc<204) then grbp<="010";
	end if;
	if (ll=218 and cc>=241 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=219) then grbp<="010";
	end if;
	if (ll=219 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=219 and cc>=28 and cc<52) then grbp<="010";
	end if;
	if (ll=219 and cc>=56 and cc<60) then grbp<="010";
	end if;
	if (ll=219 and cc>=61 and cc<66) then grbp<="010";
	end if;
	if (cc=80 and ll=219) then grbp<="010";
	end if;
	if (cc=90 and ll=219) then grbp<="010";
	end if;
	if (cc=105 and ll=219) then grbp<="010";
	end if;
	if (ll=219 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=219 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (cc=131 and ll=219) then grbp<="010";
	end if;
	if (ll=219 and cc>=131 and cc<133) then grbp<="010";
	end if;
	if (cc=139 and ll=219) then grbp<="010";
	end if;
	if (ll=219 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (cc=162 and ll=219) then grbp<="010";
	end if;
	if (cc=166 and ll=219) then grbp<="010";
	end if;
	if (cc=179 and ll=219) then grbp<="010";
	end if;
	if (cc=182 and ll=219) then grbp<="010";
	end if;
	if (ll=219 and cc>=182 and cc<184) then grbp<="010";
	end if;
	if (ll=219 and cc>=198 and cc<204) then grbp<="010";
	end if;
	if (ll=219 and cc>=239 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=220) then grbp<="010";
	end if;
	if (ll=220 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=220 and cc>=28 and cc<52) then grbp<="010";
	end if;
	if (ll=220 and cc>=55 and cc<65) then grbp<="010";
	end if;
	if (cc=118 and ll=220) then grbp<="010";
	end if;
	if (ll=220 and cc>=118 and cc<122) then grbp<="010";
	end if;
	if (ll=220 and cc>=125 and cc<127) then grbp<="010";
	end if;
	if (cc=131 and ll=220) then grbp<="010";
	end if;
	if (cc=137 and ll=220) then grbp<="010";
	end if;
	if (cc=139 and ll=220) then grbp<="010";
	end if;
	if (ll=220 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (cc=166 and ll=220) then grbp<="010";
	end if;
	if (cc=179 and ll=220) then grbp<="010";
	end if;
	if (cc=182 and ll=220) then grbp<="010";
	end if;
	if (ll=220 and cc>=182 and cc<184) then grbp<="010";
	end if;
	if (ll=220 and cc>=198 and cc<203) then grbp<="010";
	end if;
	if (ll=220 and cc>=233 and cc<235) then grbp<="010";
	end if;
	if (ll=220 and cc>=239 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=221) then grbp<="010";
	end if;
	if (ll=221 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=221 and cc>=28 and cc<53) then grbp<="010";
	end if;
	if (ll=221 and cc>=56 and cc<64) then grbp<="010";
	end if;
	if (cc=79 and ll=221) then grbp<="010";
	end if;
	if (cc=104 and ll=221) then grbp<="010";
	end if;
	if (ll=221 and cc>=104 and cc<107) then grbp<="010";
	end if;
	if (ll=221 and cc>=118 and cc<121) then grbp<="010";
	end if;
	if (ll=221 and cc>=125 and cc<127) then grbp<="010";
	end if;
	if (cc=131 and ll=221) then grbp<="010";
	end if;
	if (cc=138 and ll=221) then grbp<="010";
	end if;
	if (ll=221 and cc>=138 and cc<150) then grbp<="010";
	end if;
	if (cc=163 and ll=221) then grbp<="010";
	end if;
	if (cc=166 and ll=221) then grbp<="010";
	end if;
	if (ll=221 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=182 and ll=221) then grbp<="010";
	end if;
	if (ll=221 and cc>=182 and cc<184) then grbp<="010";
	end if;
	if (ll=221 and cc>=198 and cc<203) then grbp<="010";
	end if;
	if (ll=221 and cc>=233 and cc<235) then grbp<="010";
	end if;
	if (ll=221 and cc>=236 and cc<240) then grbp<="010";
	end if;
	if (ll=221 and cc>=241 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=222 and cc>=29 and cc<51) then grbp<="010";
	end if;
	if (cc=54 and ll=222) then grbp<="010";
	end if;
	if (cc=58 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=58 and cc<64) then grbp<="010";
	end if;
	if (cc=104 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=104 and cc<107) then grbp<="010";
	end if;
	if (ll=222 and cc>=117 and cc<122) then grbp<="010";
	end if;
	if (ll=222 and cc>=125 and cc<127) then grbp<="010";
	end if;
	if (ll=222 and cc>=128 and cc<132) then grbp<="010";
	end if;
	if (ll=222 and cc>=138 and cc<150) then grbp<="010";
	end if;
	if (ll=222 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (cc=161 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=161 and cc<163) then grbp<="010";
	end if;
	if (ll=222 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=222) then grbp<="010";
	end if;
	if (cc=182 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=182 and cc<184) then grbp<="010";
	end if;
	if (cc=197 and ll=222) then grbp<="010";
	end if;
	if (ll=222 and cc>=197 and cc<203) then grbp<="010";
	end if;
	if (ll=222 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (ll=222 and cc>=237 and cc<240) then grbp<="010";
	end if;
	if (ll=222 and cc>=241 and cc<249) then grbp<="010";
	end if;
	if (ll=223 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=223 and cc>=28 and cc<51) then grbp<="010";
	end if;
	if (cc=54 and ll=223) then grbp<="010";
	end if;
	if (ll=223 and cc>=54 and cc<56) then grbp<="010";
	end if;
	if (ll=223 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (cc=104 and ll=223) then grbp<="010";
	end if;
	if (ll=223 and cc>=104 and cc<106) then grbp<="010";
	end if;
	if (ll=223 and cc>=117 and cc<123) then grbp<="010";
	end if;
	if (ll=223 and cc>=125 and cc<128) then grbp<="010";
	end if;
	if (ll=223 and cc>=129 and cc<131) then grbp<="010";
	end if;
	if (cc=138 and ll=223) then grbp<="010";
	end if;
	if (ll=223 and cc>=138 and cc<149) then grbp<="010";
	end if;
	if (ll=223 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (ll=223 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=223 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=223) then grbp<="010";
	end if;
	if (cc=182 and ll=223) then grbp<="010";
	end if;
	if (ll=223 and cc>=182 and cc<185) then grbp<="010";
	end if;
	if (ll=223 and cc>=197 and cc<203) then grbp<="010";
	end if;
	if (cc=233 and ll=223) then grbp<="010";
	end if;
	if (ll=223 and cc>=233 and cc<249) then grbp<="010";
	end if;
	if (ll=224 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=224 and cc>=28 and cc<50) then grbp<="010";
	end if;
	if (cc=60 and ll=224) then grbp<="010";
	end if;
	if (cc=67 and ll=224) then grbp<="010";
	end if;
	if (cc=103 and ll=224) then grbp<="010";
	end if;
	if (ll=224 and cc>=103 and cc<106) then grbp<="010";
	end if;
	if (ll=224 and cc>=116 and cc<124) then grbp<="010";
	end if;
	if (ll=224 and cc>=125 and cc<128) then grbp<="010";
	end if;
	if (ll=224 and cc>=138 and cc<149) then grbp<="010";
	end if;
	if (ll=224 and cc>=155 and cc<162) then grbp<="010";
	end if;
	if (ll=224 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=224) then grbp<="010";
	end if;
	if (cc=182 and ll=224) then grbp<="010";
	end if;
	if (ll=224 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=224 and cc>=197 and cc<203) then grbp<="010";
	end if;
	if (cc=214 and ll=224) then grbp<="010";
	end if;
	if (cc=230 and ll=224) then grbp<="010";
	end if;
	if (ll=224 and cc>=230 and cc<232) then grbp<="010";
	end if;
	if (cc=235 and ll=224) then grbp<="010";
	end if;
	if (ll=224 and cc>=235 and cc<248) then grbp<="010";
	end if;
	if (ll=225 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=225 and cc>=28 and cc<49) then grbp<="010";
	end if;
	if (cc=79 and ll=225) then grbp<="010";
	end if;
	if (ll=225 and cc>=79 and cc<81) then grbp<="010";
	end if;
	if (ll=225 and cc>=103 and cc<106) then grbp<="010";
	end if;
	if (ll=225 and cc>=116 and cc<124) then grbp<="010";
	end if;
	if (ll=225 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=225 and cc>=138 and cc<149) then grbp<="010";
	end if;
	if (ll=225 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (ll=225 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=225 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=225) then grbp<="010";
	end if;
	if (cc=182 and ll=225) then grbp<="010";
	end if;
	if (cc=184 and ll=225) then grbp<="010";
	end if;
	if (ll=225 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=225 and cc>=197 and cc<202) then grbp<="010";
	end if;
	if (cc=233 and ll=225) then grbp<="010";
	end if;
	if (ll=225 and cc>=233 and cc<239) then grbp<="010";
	end if;
	if (ll=225 and cc>=240 and cc<246) then grbp<="010";
	end if;
	if (ll=226 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=226 and cc>=29 and cc<48) then grbp<="010";
	end if;
	if (ll=226 and cc>=51 and cc<53) then grbp<="010";
	end if;
	if (cc=67 and ll=226) then grbp<="010";
	end if;
	if (cc=80 and ll=226) then grbp<="010";
	end if;
	if (cc=102 and ll=226) then grbp<="010";
	end if;
	if (ll=226 and cc>=102 and cc<105) then grbp<="010";
	end if;
	if (ll=226 and cc>=115 and cc<128) then grbp<="010";
	end if;
	if (cc=137 and ll=226) then grbp<="010";
	end if;
	if (ll=226 and cc>=137 and cc<150) then grbp<="010";
	end if;
	if (ll=226 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (ll=226 and cc>=159 and cc<162) then grbp<="010";
	end if;
	if (ll=226 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=226) then grbp<="010";
	end if;
	if (cc=182 and ll=226) then grbp<="010";
	end if;
	if (cc=184 and ll=226) then grbp<="010";
	end if;
	if (ll=226 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=226 and cc>=197 and cc<202) then grbp<="010";
	end if;
	if (cc=232 and ll=226) then grbp<="010";
	end if;
	if (ll=226 and cc>=232 and cc<245) then grbp<="010";
	end if;
	if (ll=227 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=227 and cc>=29 and cc<46) then grbp<="010";
	end if;
	if (ll=227 and cc>=49 and cc<51) then grbp<="010";
	end if;
	if (cc=74 and ll=227) then grbp<="010";
	end if;
	if (cc=102 and ll=227) then grbp<="010";
	end if;
	if (ll=227 and cc>=102 and cc<105) then grbp<="010";
	end if;
	if (ll=227 and cc>=114 and cc<129) then grbp<="010";
	end if;
	if (ll=227 and cc>=138 and cc<149) then grbp<="010";
	end if;
	if (ll=227 and cc>=155 and cc<159) then grbp<="010";
	end if;
	if (ll=227 and cc>=165 and cc<168) then grbp<="010";
	end if;
	if (cc=179 and ll=227) then grbp<="010";
	end if;
	if (cc=182 and ll=227) then grbp<="010";
	end if;
	if (cc=184 and ll=227) then grbp<="010";
	end if;
	if (cc=197 and ll=227) then grbp<="010";
	end if;
	if (ll=227 and cc>=197 and cc<202) then grbp<="010";
	end if;
	if (cc=228 and ll=227) then grbp<="010";
	end if;
	if (ll=227 and cc>=228 and cc<232) then grbp<="010";
	end if;
	if (ll=227 and cc>=233 and cc<243) then grbp<="010";
	end if;
	if (ll=228 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=228 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=57 and ll=228) then grbp<="010";
	end if;
	if (cc=67 and ll=228) then grbp<="010";
	end if;
	if (cc=102 and ll=228) then grbp<="010";
	end if;
	if (ll=228 and cc>=102 and cc<105) then grbp<="010";
	end if;
	if (ll=228 and cc>=114 and cc<130) then grbp<="010";
	end if;
	if (ll=228 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=228 and cc>=156 and cc<159) then grbp<="010";
	end if;
	if (ll=228 and cc>=164 and cc<167) then grbp<="010";
	end if;
	if (cc=177 and ll=228) then grbp<="010";
	end if;
	if (cc=182 and ll=228) then grbp<="010";
	end if;
	if (ll=228 and cc>=182 and cc<185) then grbp<="010";
	end if;
	if (ll=228 and cc>=196 and cc<202) then grbp<="010";
	end if;
	if (cc=228 and ll=228) then grbp<="010";
	end if;
	if (ll=228 and cc>=228 and cc<243) then grbp<="010";
	end if;
	if (ll=229 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=229 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=101 and ll=229) then grbp<="010";
	end if;
	if (ll=229 and cc>=101 and cc<104) then grbp<="010";
	end if;
	if (ll=229 and cc>=113 and cc<134) then grbp<="010";
	end if;
	if (ll=229 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=229 and cc>=158 and cc<162) then grbp<="010";
	end if;
	if (ll=229 and cc>=164 and cc<167) then grbp<="010";
	end if;
	if (cc=177 and ll=229) then grbp<="010";
	end if;
	if (cc=182 and ll=229) then grbp<="010";
	end if;
	if (ll=229 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=229 and cc>=196 and cc<202) then grbp<="010";
	end if;
	if (ll=229 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (cc=226 and ll=229) then grbp<="010";
	end if;
	if (ll=229 and cc>=226 and cc<228) then grbp<="010";
	end if;
	if (ll=229 and cc>=229 and cc<242) then grbp<="010";
	end if;
	if (ll=230 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=230 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (ll=230 and cc>=47 and cc<49) then grbp<="010";
	end if;
	if (cc=101 and ll=230) then grbp<="010";
	end if;
	if (ll=230 and cc>=101 and cc<104) then grbp<="010";
	end if;
	if (ll=230 and cc>=112 and cc<136) then grbp<="010";
	end if;
	if (ll=230 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=230 and cc>=157 and cc<171) then grbp<="010";
	end if;
	if (cc=183 and ll=230) then grbp<="010";
	end if;
	if (ll=230 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=230 and cc>=196 and cc<202) then grbp<="010";
	end if;
	if (cc=226 and ll=230) then grbp<="010";
	end if;
	if (ll=230 and cc>=226 and cc<240) then grbp<="010";
	end if;
	if (ll=231 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=231 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (ll=231 and cc>=47 and cc<49) then grbp<="010";
	end if;
	if (cc=63 and ll=231) then grbp<="010";
	end if;
	if (cc=101 and ll=231) then grbp<="010";
	end if;
	if (ll=231 and cc>=101 and cc<104) then grbp<="010";
	end if;
	if (ll=231 and cc>=112 and cc<134) then grbp<="010";
	end if;
	if (cc=139 and ll=231) then grbp<="010";
	end if;
	if (ll=231 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (ll=231 and cc>=156 and cc<171) then grbp<="010";
	end if;
	if (cc=183 and ll=231) then grbp<="010";
	end if;
	if (ll=231 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=231 and cc>=196 and cc<201) then grbp<="010";
	end if;
	if (ll=231 and cc>=226 and cc<239) then grbp<="010";
	end if;
	if (ll=232 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=232 and cc>=29 and cc<49) then grbp<="010";
	end if;
	if (ll=232 and cc>=52 and cc<56) then grbp<="010";
	end if;
	if (ll=232 and cc>=100 and cc<104) then grbp<="010";
	end if;
	if (ll=232 and cc>=111 and cc<134) then grbp<="010";
	end if;
	if (cc=139 and ll=232) then grbp<="010";
	end if;
	if (ll=232 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (ll=232 and cc>=156 and cc<171) then grbp<="010";
	end if;
	if (ll=232 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (ll=232 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (cc=227 and ll=232) then grbp<="010";
	end if;
	if (ll=232 and cc>=227 and cc<238) then grbp<="010";
	end if;
	if (ll=233 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=233 and cc>=29 and cc<46) then grbp<="010";
	end if;
	if (cc=55 and ll=233) then grbp<="010";
	end if;
	if (cc=100 and ll=233) then grbp<="010";
	end if;
	if (ll=233 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=233 and cc>=111 and cc<135) then grbp<="010";
	end if;
	if (ll=233 and cc>=141 and cc<150) then grbp<="010";
	end if;
	if (ll=233 and cc>=158 and cc<171) then grbp<="010";
	end if;
	if (cc=195 and ll=233) then grbp<="010";
	end if;
	if (ll=233 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (cc=225 and ll=233) then grbp<="010";
	end if;
	if (ll=233 and cc>=225 and cc<238) then grbp<="010";
	end if;
	if (ll=234 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=234 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=50 and ll=234) then grbp<="010";
	end if;
	if (ll=234 and cc>=50 and cc<52) then grbp<="010";
	end if;
	if (cc=63 and ll=234) then grbp<="010";
	end if;
	if (cc=100 and ll=234) then grbp<="010";
	end if;
	if (ll=234 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=234 and cc>=110 and cc<120) then grbp<="010";
	end if;
	if (ll=234 and cc>=121 and cc<133) then grbp<="010";
	end if;
	if (ll=234 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=234 and cc>=158 and cc<171) then grbp<="010";
	end if;
	if (cc=195 and ll=234) then grbp<="010";
	end if;
	if (ll=234 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (cc=214 and ll=234) then grbp<="010";
	end if;
	if (cc=224 and ll=234) then grbp<="010";
	end if;
	if (ll=234 and cc>=224 and cc<237) then grbp<="010";
	end if;
	if (ll=235 and cc>=0 and cc<12) then grbp<="010";
	end if;
	if (ll=235 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=235 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (ll=235 and cc>=49 and cc<51) then grbp<="010";
	end if;
	if (cc=80 and ll=235) then grbp<="010";
	end if;
	if (cc=99 and ll=235) then grbp<="010";
	end if;
	if (ll=235 and cc>=99 and cc<103) then grbp<="010";
	end if;
	if (ll=235 and cc>=110 and cc<118) then grbp<="010";
	end if;
	if (ll=235 and cc>=119 and cc<123) then grbp<="010";
	end if;
	if (ll=235 and cc>=124 and cc<133) then grbp<="010";
	end if;
	if (ll=235 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=235 and cc>=159 and cc<171) then grbp<="010";
	end if;
	if (cc=195 and ll=235) then grbp<="010";
	end if;
	if (ll=235 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (cc=224 and ll=235) then grbp<="010";
	end if;
	if (ll=235 and cc>=224 and cc<236) then grbp<="010";
	end if;
	if (ll=236 and cc>=0 and cc<12) then grbp<="010";
	end if;
	if (ll=236 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=236 and cc>=29 and cc<46) then grbp<="010";
	end if;
	if (ll=236 and cc>=48 and cc<51) then grbp<="010";
	end if;
	if (cc=67 and ll=236) then grbp<="010";
	end if;
	if (cc=99 and ll=236) then grbp<="010";
	end if;
	if (ll=236 and cc>=99 and cc<102) then grbp<="010";
	end if;
	if (ll=236 and cc>=109 and cc<121) then grbp<="010";
	end if;
	if (ll=236 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=236 and cc>=160 and cc<172) then grbp<="010";
	end if;
	if (cc=185 and ll=236) then grbp<="010";
	end if;
	if (cc=195 and ll=236) then grbp<="010";
	end if;
	if (ll=236 and cc>=195 and cc<201) then grbp<="010";
	end if;
	if (ll=236 and cc>=223 and cc<235) then grbp<="010";
	end if;
	if (ll=237 and cc>=0 and cc<12) then grbp<="010";
	end if;
	if (ll=237 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=237 and cc>=29 and cc<51) then grbp<="010";
	end if;
	if (cc=67 and ll=237) then grbp<="010";
	end if;
	if (cc=99 and ll=237) then grbp<="010";
	end if;
	if (ll=237 and cc>=99 and cc<102) then grbp<="010";
	end if;
	if (ll=237 and cc>=109 and cc<120) then grbp<="010";
	end if;
	if (ll=237 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=237 and cc>=160 and cc<172) then grbp<="010";
	end if;
	if (cc=185 and ll=237) then grbp<="010";
	end if;
	if (cc=195 and ll=237) then grbp<="010";
	end if;
	if (ll=237 and cc>=195 and cc<200) then grbp<="010";
	end if;
	if (cc=217 and ll=237) then grbp<="010";
	end if;
	if (cc=220 and ll=237) then grbp<="010";
	end if;
	if (ll=237 and cc>=220 and cc<235) then grbp<="010";
	end if;
	if (ll=238 and cc>=0 and cc<12) then grbp<="010";
	end if;
	if (ll=238 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=238 and cc>=29 and cc<50) then grbp<="010";
	end if;
	if (cc=83 and ll=238) then grbp<="010";
	end if;
	if (cc=98 and ll=238) then grbp<="010";
	end if;
	if (ll=238 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=238 and cc>=108 and cc<120) then grbp<="010";
	end if;
	if (ll=238 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=238 and cc>=160 and cc<172) then grbp<="010";
	end if;
	if (cc=185 and ll=238) then grbp<="010";
	end if;
	if (cc=195 and ll=238) then grbp<="010";
	end if;
	if (ll=238 and cc>=195 and cc<200) then grbp<="010";
	end if;
	if (ll=238 and cc>=209 and cc<211) then grbp<="010";
	end if;
	if (cc=222 and ll=238) then grbp<="010";
	end if;
	if (cc=224 and ll=238) then grbp<="010";
	end if;
	if (ll=238 and cc>=224 and cc<234) then grbp<="010";
	end if;
	if (ll=239 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=239 and cc>=29 and cc<47) then grbp<="010";
	end if;
	if (cc=74 and ll=239) then grbp<="010";
	end if;
	if (cc=98 and ll=239) then grbp<="010";
	end if;
	if (ll=239 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=239 and cc>=109 and cc<120) then grbp<="010";
	end if;
	if (ll=239 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (ll=239 and cc>=160 and cc<171) then grbp<="010";
	end if;
	if (cc=183 and ll=239) then grbp<="010";
	end if;
	if (cc=185 and ll=239) then grbp<="010";
	end if;
	if (cc=194 and ll=239) then grbp<="010";
	end if;
	if (ll=239 and cc>=194 and cc<200) then grbp<="010";
	end if;
	if (ll=239 and cc>=207 and cc<210) then grbp<="010";
	end if;
	if (cc=221 and ll=239) then grbp<="010";
	end if;
	if (ll=239 and cc>=221 and cc<234) then grbp<="010";
	end if;
	if (ll=240 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=240 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=240 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=66 and ll=240) then grbp<="010";
	end if;
	if (cc=99 and ll=240) then grbp<="010";
	end if;
	if (ll=240 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (cc=109 and ll=240) then grbp<="010";
	end if;
	if (ll=240 and cc>=109 and cc<119) then grbp<="010";
	end if;
	if (ll=240 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (ll=240 and cc>=160 and cc<171) then grbp<="010";
	end if;
	if (cc=194 and ll=240) then grbp<="010";
	end if;
	if (ll=240 and cc>=194 and cc<200) then grbp<="010";
	end if;
	if (ll=240 and cc>=219 and cc<233) then grbp<="010";
	end if;
	if (ll=241 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=241 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=241 and cc>=29 and cc<42) then grbp<="010";
	end if;
	if (cc=83 and ll=241) then grbp<="010";
	end if;
	if (ll=241 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=241 and cc>=97 and cc<101) then grbp<="010";
	end if;
	if (ll=241 and cc>=108 and cc<121) then grbp<="010";
	end if;
	if (ll=241 and cc>=139 and cc<150) then grbp<="010";
	end if;
	if (ll=241 and cc>=160 and cc<171) then grbp<="010";
	end if;
	if (cc=194 and ll=241) then grbp<="010";
	end if;
	if (ll=241 and cc>=194 and cc<199) then grbp<="010";
	end if;
	if (ll=241 and cc>=219 and cc<232) then grbp<="010";
	end if;
	if (ll=242 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=242 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=242 and cc>=29 and cc<41) then grbp<="010";
	end if;
	if (cc=83 and ll=242) then grbp<="010";
	end if;
	if (ll=242 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=242 and cc>=97 and cc<101) then grbp<="010";
	end if;
	if (cc=108 and ll=242) then grbp<="010";
	end if;
	if (ll=242 and cc>=108 and cc<121) then grbp<="010";
	end if;
	if (ll=242 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (ll=242 and cc>=161 and cc<171) then grbp<="010";
	end if;
	if (ll=242 and cc>=194 and cc<199) then grbp<="010";
	end if;
	if (cc=220 and ll=242) then grbp<="010";
	end if;
	if (ll=242 and cc>=220 and cc<222) then grbp<="010";
	end if;
	if (ll=242 and cc>=223 and cc<232) then grbp<="010";
	end if;
	if (ll=243 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=243 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=243 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (cc=46 and ll=243) then grbp<="010";
	end if;
	if (ll=243 and cc>=46 and cc<48) then grbp<="010";
	end if;
	if (cc=85 and ll=243) then grbp<="010";
	end if;
	if (ll=243 and cc>=85 and cc<87) then grbp<="010";
	end if;
	if (ll=243 and cc>=98 and cc<100) then grbp<="010";
	end if;
	if (ll=243 and cc>=108 and cc<121) then grbp<="010";
	end if;
	if (ll=243 and cc>=140 and cc<151) then grbp<="010";
	end if;
	if (ll=243 and cc>=160 and cc<171) then grbp<="010";
	end if;
	if (cc=194 and ll=243) then grbp<="010";
	end if;
	if (ll=243 and cc>=194 and cc<199) then grbp<="010";
	end if;
	if (ll=243 and cc>=212 and cc<214) then grbp<="010";
	end if;
	if (ll=243 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=243 and cc>=220 and cc<232) then grbp<="010";
	end if;
	if (ll=244 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=244 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=244 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (ll=244 and cc>=40 and cc<43) then grbp<="010";
	end if;
	if (ll=244 and cc>=46 and cc<48) then grbp<="010";
	end if;
	if (cc=83 and ll=244) then grbp<="010";
	end if;
	if (ll=244 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=244 and cc>=97 and cc<100) then grbp<="010";
	end if;
	if (ll=244 and cc>=108 and cc<122) then grbp<="010";
	end if;
	if (ll=244 and cc>=140 and cc<150) then grbp<="010";
	end if;
	if (ll=244 and cc>=160 and cc<171) then grbp<="010";
	end if;
	if (cc=194 and ll=244) then grbp<="010";
	end if;
	if (ll=244 and cc>=194 and cc<199) then grbp<="010";
	end if;
	if (ll=244 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=244 and cc>=222 and cc<231) then grbp<="010";
	end if;
	if (ll=245 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=245 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=245 and cc>=29 and cc<43) then grbp<="010";
	end if;
	if (cc=47 and ll=245) then grbp<="010";
	end if;
	if (cc=78 and ll=245) then grbp<="010";
	end if;
	if (cc=82 and ll=245) then grbp<="010";
	end if;
	if (ll=245 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=245 and cc>=96 and cc<100) then grbp<="010";
	end if;
	if (ll=245 and cc>=108 and cc<122) then grbp<="010";
	end if;
	if (ll=245 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (ll=245 and cc>=161 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=245) then grbp<="010";
	end if;
	if (cc=182 and ll=245) then grbp<="010";
	end if;
	if (cc=193 and ll=245) then grbp<="010";
	end if;
	if (ll=245 and cc>=193 and cc<199) then grbp<="010";
	end if;
	if (cc=217 and ll=245) then grbp<="010";
	end if;
	if (cc=219 and ll=245) then grbp<="010";
	end if;
	if (cc=221 and ll=245) then grbp<="010";
	end if;
	if (ll=245 and cc>=221 and cc<231) then grbp<="010";
	end if;
	if (ll=246 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=246 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=246 and cc>=29 and cc<50) then grbp<="010";
	end if;
	if (cc=82 and ll=246) then grbp<="010";
	end if;
	if (ll=246 and cc>=82 and cc<87) then grbp<="010";
	end if;
	if (ll=246 and cc>=96 and cc<99) then grbp<="010";
	end if;
	if (ll=246 and cc>=108 and cc<122) then grbp<="010";
	end if;
	if (ll=246 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (ll=246 and cc>=161 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=246) then grbp<="010";
	end if;
	if (cc=182 and ll=246) then grbp<="010";
	end if;
	if (cc=184 and ll=246) then grbp<="010";
	end if;
	if (cc=193 and ll=246) then grbp<="010";
	end if;
	if (ll=246 and cc>=193 and cc<198) then grbp<="010";
	end if;
	if (cc=213 and ll=246) then grbp<="010";
	end if;
	if (ll=246 and cc>=213 and cc<216) then grbp<="010";
	end if;
	if (ll=246 and cc>=219 and cc<221) then grbp<="010";
	end if;
	if (ll=246 and cc>=222 and cc<231) then grbp<="010";
	end if;
	if (ll=247 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=247 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=247 and cc>=28 and cc<46) then grbp<="010";
	end if;
	if (cc=61 and ll=247) then grbp<="010";
	end if;
	if (cc=83 and ll=247) then grbp<="010";
	end if;
	if (ll=247 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=247 and cc>=97 and cc<99) then grbp<="010";
	end if;
	if (cc=108 and ll=247) then grbp<="010";
	end if;
	if (ll=247 and cc>=108 and cc<122) then grbp<="010";
	end if;
	if (ll=247 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=247 and cc>=161 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=247) then grbp<="010";
	end if;
	if (cc=182 and ll=247) then grbp<="010";
	end if;
	if (cc=184 and ll=247) then grbp<="010";
	end if;
	if (cc=193 and ll=247) then grbp<="010";
	end if;
	if (ll=247 and cc>=193 and cc<198) then grbp<="010";
	end if;
	if (cc=213 and ll=247) then grbp<="010";
	end if;
	if (ll=247 and cc>=213 and cc<216) then grbp<="010";
	end if;
	if (cc=219 and ll=247) then grbp<="010";
	end if;
	if (cc=221 and ll=247) then grbp<="010";
	end if;
	if (ll=247 and cc>=221 and cc<230) then grbp<="010";
	end if;
	if (ll=248 and cc>=0 and cc<10) then grbp<="010";
	end if;
	if (ll=248 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=248 and cc>=28 and cc<46) then grbp<="010";
	end if;
	if (cc=83 and ll=248) then grbp<="010";
	end if;
	if (ll=248 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=248 and cc>=95 and cc<99) then grbp<="010";
	end if;
	if (ll=248 and cc>=108 and cc<123) then grbp<="010";
	end if;
	if (ll=248 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=248 and cc>=161 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=248) then grbp<="010";
	end if;
	if (cc=182 and ll=248) then grbp<="010";
	end if;
	if (cc=184 and ll=248) then grbp<="010";
	end if;
	if (cc=193 and ll=248) then grbp<="010";
	end if;
	if (ll=248 and cc>=193 and cc<198) then grbp<="010";
	end if;
	if (cc=211 and ll=248) then grbp<="010";
	end if;
	if (cc=215 and ll=248) then grbp<="010";
	end if;
	if (cc=217 and ll=248) then grbp<="010";
	end if;
	if (cc=219 and ll=248) then grbp<="010";
	end if;
	if (ll=248 and cc>=219 and cc<230) then grbp<="010";
	end if;
	if (ll=249 and cc>=0 and cc<10) then grbp<="010";
	end if;
	if (ll=249 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=249 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (ll=249 and cc>=50 and cc<52) then grbp<="010";
	end if;
	if (ll=249 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (cc=95 and ll=249) then grbp<="010";
	end if;
	if (ll=249 and cc>=95 and cc<99) then grbp<="010";
	end if;
	if (cc=108 and ll=249) then grbp<="010";
	end if;
	if (ll=249 and cc>=108 and cc<123) then grbp<="010";
	end if;
	if (ll=249 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=249 and cc>=162 and cc<171) then grbp<="010";
	end if;
	if (cc=180 and ll=249) then grbp<="010";
	end if;
	if (cc=184 and ll=249) then grbp<="010";
	end if;
	if (cc=193 and ll=249) then grbp<="010";
	end if;
	if (ll=249 and cc>=193 and cc<197) then grbp<="010";
	end if;
	if (ll=249 and cc>=213 and cc<215) then grbp<="010";
	end if;
	if (ll=249 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=249 and cc>=220 and cc<229) then grbp<="010";
	end if;
	if (ll=250 and cc>=0 and cc<10) then grbp<="010";
	end if;
	if (ll=250 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=250 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=50 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=50 and cc<52) then grbp<="010";
	end if;
	if (cc=82 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (cc=95 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=95 and cc<98) then grbp<="010";
	end if;
	if (ll=250 and cc>=108 and cc<124) then grbp<="010";
	end if;
	if (ll=250 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (ll=250 and cc>=160 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=250) then grbp<="010";
	end if;
	if (cc=193 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=193 and cc<197) then grbp<="010";
	end if;
	if (cc=213 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=213 and cc<229) then grbp<="010";
	end if;
	if (ll=251 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (cc=13 and ll=251) then grbp<="010";
	end if;
	if (ll=251 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=251 and cc>=29 and cc<44) then grbp<="010";
	end if;
	if (cc=49 and ll=251) then grbp<="010";
	end if;
	if (cc=51 and ll=251) then grbp<="010";
	end if;
	if (cc=82 and ll=251) then grbp<="010";
	end if;
	if (ll=251 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (cc=94 and ll=251) then grbp<="010";
	end if;
	if (ll=251 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=251 and cc>=108 and cc<124) then grbp<="010";
	end if;
	if (ll=251 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=251 and cc>=160 and cc<162) then grbp<="010";
	end if;
	if (ll=251 and cc>=163 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=251) then grbp<="010";
	end if;
	if (cc=192 and ll=251) then grbp<="010";
	end if;
	if (ll=251 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (ll=251 and cc>=209 and cc<211) then grbp<="010";
	end if;
	if (ll=251 and cc>=212 and cc<215) then grbp<="010";
	end if;
	if (ll=251 and cc>=216 and cc<229) then grbp<="010";
	end if;
	if (ll=252 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=252 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=252 and cc>=28 and cc<36) then grbp<="010";
	end if;
	if (ll=252 and cc>=37 and cc<43) then grbp<="010";
	end if;
	if (cc=82 and ll=252) then grbp<="010";
	end if;
	if (ll=252 and cc>=82 and cc<89) then grbp<="010";
	end if;
	if (ll=252 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (cc=108 and ll=252) then grbp<="010";
	end if;
	if (ll=252 and cc>=108 and cc<125) then grbp<="010";
	end if;
	if (ll=252 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=252 and cc>=160 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=252) then grbp<="010";
	end if;
	if (cc=192 and ll=252) then grbp<="010";
	end if;
	if (ll=252 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (cc=212 and ll=252) then grbp<="010";
	end if;
	if (ll=252 and cc>=212 and cc<218) then grbp<="010";
	end if;
	if (ll=252 and cc>=219 and cc<228) then grbp<="010";
	end if;
	if (ll=253 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=253 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=253 and cc>=28 and cc<36) then grbp<="010";
	end if;
	if (ll=253 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=82 and ll=253) then grbp<="010";
	end if;
	if (cc=84 and ll=253) then grbp<="010";
	end if;
	if (ll=253 and cc>=84 and cc<88) then grbp<="010";
	end if;
	if (cc=94 and ll=253) then grbp<="010";
	end if;
	if (ll=253 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=253 and cc>=108 and cc<125) then grbp<="010";
	end if;
	if (ll=253 and cc>=137 and cc<151) then grbp<="010";
	end if;
	if (ll=253 and cc>=160 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=253) then grbp<="010";
	end if;
	if (cc=184 and ll=253) then grbp<="010";
	end if;
	if (cc=192 and ll=253) then grbp<="010";
	end if;
	if (ll=253 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (ll=253 and cc>=210 and cc<228) then grbp<="010";
	end if;
	if (ll=254 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=254 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=254 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=254 and cc>=37 and cc<40) then grbp<="010";
	end if;
	if (cc=50 and ll=254) then grbp<="010";
	end if;
	if (cc=52 and ll=254) then grbp<="010";
	end if;
	if (cc=62 and ll=254) then grbp<="010";
	end if;
	if (cc=76 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=254 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (cc=87 and ll=254) then grbp<="010";
	end if;
	if (cc=89 and ll=254) then grbp<="010";
	end if;
	if (cc=94 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=254 and cc>=108 and cc<123) then grbp<="010";
	end if;
	if (cc=138 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=138 and cc<151) then grbp<="010";
	end if;
	if (ll=254 and cc>=160 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=254) then grbp<="010";
	end if;
	if (cc=185 and ll=254) then grbp<="010";
	end if;
	if (cc=192 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (cc=214 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=214 and cc<228) then grbp<="010";
	end if;
	if (ll=255 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=255 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=255 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=255 and cc>=37 and cc<39) then grbp<="010";
	end if;
	if (cc=44 and ll=255) then grbp<="010";
	end if;
	if (cc=47 and ll=255) then grbp<="010";
	end if;
	if (cc=50 and ll=255) then grbp<="010";
	end if;
	if (cc=76 and ll=255) then grbp<="010";
	end if;
	if (ll=255 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=255 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (cc=87 and ll=255) then grbp<="010";
	end if;
	if (ll=255 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=255 and cc>=93 and cc<97) then grbp<="010";
	end if;
	if (cc=108 and ll=255) then grbp<="010";
	end if;
	if (ll=255 and cc>=108 and cc<125) then grbp<="010";
	end if;
	if (ll=255 and cc>=137 and cc<151) then grbp<="010";
	end if;
	if (ll=255 and cc>=161 and cc<170) then grbp<="010";
	end if;
	if (cc=180 and ll=255) then grbp<="010";
	end if;
	if (cc=184 and ll=255) then grbp<="010";
	end if;
	if (ll=255 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=255 and cc>=192 and cc<197) then grbp<="010";
	end if;
	if (ll=255 and cc>=212 and cc<214) then grbp<="010";
	end if;
	if (ll=255 and cc>=216 and cc<227) then grbp<="010";
	end if;
	if (ll=256 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=256 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=256 and cc>=29 and cc<37) then grbp<="010";
	end if;
	if (cc=41 and ll=256) then grbp<="010";
	end if;
	if (cc=44 and ll=256) then grbp<="010";
	end if;
	if (cc=49 and ll=256) then grbp<="010";
	end if;
	if (cc=76 and ll=256) then grbp<="010";
	end if;
	if (ll=256 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (cc=85 and ll=256) then grbp<="010";
	end if;
	if (cc=87 and ll=256) then grbp<="010";
	end if;
	if (ll=256 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=256 and cc>=93 and cc<97) then grbp<="010";
	end if;
	if (cc=108 and ll=256) then grbp<="010";
	end if;
	if (ll=256 and cc>=108 and cc<124) then grbp<="010";
	end if;
	if (ll=256 and cc>=137 and cc<151) then grbp<="010";
	end if;
	if (ll=256 and cc>=159 and cc<170) then grbp<="010";
	end if;
	if (cc=183 and ll=256) then grbp<="010";
	end if;
	if (ll=256 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=256 and cc>=192 and cc<196) then grbp<="010";
	end if;
	if (cc=212 and ll=256) then grbp<="010";
	end if;
	if (ll=256 and cc>=212 and cc<214) then grbp<="010";
	end if;
	if (ll=256 and cc>=216 and cc<227) then grbp<="010";
	end if;
	if (ll=257 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=257 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=257 and cc>=29 and cc<37) then grbp<="010";
	end if;
	if (ll=257 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=257 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (cc=50 and ll=257) then grbp<="010";
	end if;
	if (cc=76 and ll=257) then grbp<="010";
	end if;
	if (ll=257 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=257 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (cc=93 and ll=257) then grbp<="010";
	end if;
	if (ll=257 and cc>=93 and cc<97) then grbp<="010";
	end if;
	if (cc=106 and ll=257) then grbp<="010";
	end if;
	if (cc=108 and ll=257) then grbp<="010";
	end if;
	if (ll=257 and cc>=108 and cc<125) then grbp<="010";
	end if;
	if (ll=257 and cc>=137 and cc<151) then grbp<="010";
	end if;
	if (ll=257 and cc>=160 and cc<170) then grbp<="010";
	end if;
	if (cc=183 and ll=257) then grbp<="010";
	end if;
	if (ll=257 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=257 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (cc=211 and ll=257) then grbp<="010";
	end if;
	if (ll=257 and cc>=211 and cc<214) then grbp<="010";
	end if;
	if (ll=257 and cc>=216 and cc<227) then grbp<="010";
	end if;
	if (ll=258 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=258 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=258 and cc>=29 and cc<38) then grbp<="010";
	end if;
	if (ll=258 and cc>=40 and cc<45) then grbp<="010";
	end if;
	if (cc=48 and ll=258) then grbp<="010";
	end if;
	if (cc=50 and ll=258) then grbp<="010";
	end if;
	if (cc=76 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=258 and cc>=80 and cc<84) then grbp<="010";
	end if;
	if (cc=93 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (cc=108 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=108 and cc<126) then grbp<="010";
	end if;
	if (cc=137 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=137 and cc<152) then grbp<="010";
	end if;
	if (cc=159 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=159 and cc<169) then grbp<="010";
	end if;
	if (cc=183 and ll=258) then grbp<="010";
	end if;
	if (cc=185 and ll=258) then grbp<="010";
	end if;
	if (cc=191 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (cc=212 and ll=258) then grbp<="010";
	end if;
	if (cc=215 and ll=258) then grbp<="010";
	end if;
	if (ll=258 and cc>=215 and cc<218) then grbp<="010";
	end if;
	if (ll=258 and cc>=219 and cc<227) then grbp<="010";
	end if;
	if (ll=259 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=259 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=259 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (cc=48 and ll=259) then grbp<="010";
	end if;
	if (cc=77 and ll=259) then grbp<="010";
	end if;
	if (ll=259 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=259 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (cc=92 and ll=259) then grbp<="010";
	end if;
	if (ll=259 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (cc=106 and ll=259) then grbp<="010";
	end if;
	if (ll=259 and cc>=106 and cc<129) then grbp<="010";
	end if;
	if (ll=259 and cc>=137 and cc<152) then grbp<="010";
	end if;
	if (ll=259 and cc>=159 and cc<169) then grbp<="010";
	end if;
	if (cc=181 and ll=259) then grbp<="010";
	end if;
	if (cc=183 and ll=259) then grbp<="010";
	end if;
	if (ll=259 and cc>=183 and cc<186) then grbp<="010";
	end if;
	if (ll=259 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (ll=259 and cc>=215 and cc<226) then grbp<="010";
	end if;
	if (ll=260 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=260 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=260 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (cc=44 and ll=260) then grbp<="010";
	end if;
	if (cc=47 and ll=260) then grbp<="010";
	end if;
	if (cc=50 and ll=260) then grbp<="010";
	end if;
	if (cc=75 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=75 and cc<83) then grbp<="010";
	end if;
	if (cc=92 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (cc=108 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=108 and cc<129) then grbp<="010";
	end if;
	if (ll=260 and cc>=136 and cc<152) then grbp<="010";
	end if;
	if (ll=260 and cc>=158 and cc<169) then grbp<="010";
	end if;
	if (cc=181 and ll=260) then grbp<="010";
	end if;
	if (cc=183 and ll=260) then grbp<="010";
	end if;
	if (cc=185 and ll=260) then grbp<="010";
	end if;
	if (cc=191 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (ll=260 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (cc=216 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=216 and cc<226) then grbp<="010";
	end if;
	if (ll=261 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=261 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=261 and cc>=29 and cc<44) then grbp<="010";
	end if;
	if (cc=50 and ll=261) then grbp<="010";
	end if;
	if (cc=77 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=77 and cc<85) then grbp<="010";
	end if;
	if (ll=261 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (cc=108 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=108 and cc<128) then grbp<="010";
	end if;
	if (ll=261 and cc>=136 and cc<152) then grbp<="010";
	end if;
	if (ll=261 and cc>=158 and cc<169) then grbp<="010";
	end if;
	if (cc=181 and ll=261) then grbp<="010";
	end if;
	if (cc=185 and ll=261) then grbp<="010";
	end if;
	if (cc=191 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=191 and cc<196) then grbp<="010";
	end if;
	if (cc=211 and ll=261) then grbp<="010";
	end if;
	if (cc=214 and ll=261) then grbp<="010";
	end if;
	if (cc=217 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=217 and cc<225) then grbp<="010";
	end if;
	if (ll=262 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=262 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=262 and cc>=29 and cc<37) then grbp<="010";
	end if;
	if (ll=262 and cc>=39 and cc<44) then grbp<="010";
	end if;
	if (cc=50 and ll=262) then grbp<="010";
	end if;
	if (cc=65 and ll=262) then grbp<="010";
	end if;
	if (cc=77 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=77 and cc<79) then grbp<="010";
	end if;
	if (ll=262 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (ll=262 and cc>=91 and cc<95) then grbp<="010";
	end if;
	if (cc=106 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=106 and cc<130) then grbp<="010";
	end if;
	if (ll=262 and cc>=135 and cc<152) then grbp<="010";
	end if;
	if (ll=262 and cc>=158 and cc<168) then grbp<="010";
	end if;
	if (cc=181 and ll=262) then grbp<="010";
	end if;
	if (cc=185 and ll=262) then grbp<="010";
	end if;
	if (cc=190 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=190 and cc<196) then grbp<="010";
	end if;
	if (cc=217 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=217 and cc<225) then grbp<="010";
	end if;
	if (ll=263 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=263 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=263 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=263 and cc>=38 and cc<44) then grbp<="010";
	end if;
	if (ll=263 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=78 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=78 and cc<81) then grbp<="010";
	end if;
	if (cc=92 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=92 and cc<97) then grbp<="010";
	end if;
	if (cc=106 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=106 and cc<128) then grbp<="010";
	end if;
	if (ll=263 and cc>=129 and cc<131) then grbp<="010";
	end if;
	if (ll=263 and cc>=135 and cc<152) then grbp<="010";
	end if;
	if (ll=263 and cc>=158 and cc<168) then grbp<="010";
	end if;
	if (cc=181 and ll=263) then grbp<="010";
	end if;
	if (cc=185 and ll=263) then grbp<="010";
	end if;
	if (cc=190 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=190 and cc<196) then grbp<="010";
	end if;
	if (cc=213 and ll=263) then grbp<="010";
	end if;
	if (cc=218 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=218 and cc<225) then grbp<="010";
	end if;
	if (ll=264 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=264 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=264 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=264 and cc>=37 and cc<44) then grbp<="010";
	end if;
	if (cc=63 and ll=264) then grbp<="010";
	end if;
	if (cc=76 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=264 and cc>=80 and cc<83) then grbp<="010";
	end if;
	if (cc=98 and ll=264) then grbp<="010";
	end if;
	if (cc=106 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=106 and cc<127) then grbp<="010";
	end if;
	if (ll=264 and cc>=128 and cc<130) then grbp<="010";
	end if;
	if (ll=264 and cc>=136 and cc<152) then grbp<="010";
	end if;
	if (ll=264 and cc>=158 and cc<168) then grbp<="010";
	end if;
	if (ll=264 and cc>=175 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=264 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (ll=264 and cc>=209 and cc<211) then grbp<="010";
	end if;
	if (cc=216 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=216 and cc<225) then grbp<="010";
	end if;
	if (ll=265 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=265 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=265 and cc>=29 and cc<35) then grbp<="010";
	end if;
	if (ll=265 and cc>=36 and cc<44) then grbp<="010";
	end if;
	if (cc=49 and ll=265) then grbp<="010";
	end if;
	if (cc=76 and ll=265) then grbp<="010";
	end if;
	if (cc=82 and ll=265) then grbp<="010";
	end if;
	if (cc=98 and ll=265) then grbp<="010";
	end if;
	if (cc=106 and ll=265) then grbp<="010";
	end if;
	if (ll=265 and cc>=106 and cc<132) then grbp<="010";
	end if;
	if (ll=265 and cc>=134 and cc<152) then grbp<="010";
	end if;
	if (ll=265 and cc>=157 and cc<168) then grbp<="010";
	end if;
	if (cc=181 and ll=265) then grbp<="010";
	end if;
	if (cc=184 and ll=265) then grbp<="010";
	end if;
	if (ll=265 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=265 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (cc=216 and ll=265) then grbp<="010";
	end if;
	if (ll=265 and cc>=216 and cc<225) then grbp<="010";
	end if;
	if (ll=266 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=266 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=266 and cc>=29 and cc<44) then grbp<="010";
	end if;
	if (cc=81 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (cc=97 and ll=266) then grbp<="010";
	end if;
	if (cc=105 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=105 and cc<130) then grbp<="010";
	end if;
	if (cc=135 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=135 and cc<153) then grbp<="010";
	end if;
	if (ll=266 and cc>=157 and cc<167) then grbp<="010";
	end if;
	if (cc=181 and ll=266) then grbp<="010";
	end if;
	if (cc=184 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=266 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (cc=211 and ll=266) then grbp<="010";
	end if;
	if (cc=214 and ll=266) then grbp<="010";
	end if;
	if (cc=216 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=216 and cc<224) then grbp<="010";
	end if;
	if (ll=267 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=267 and cc>=13 and cc<17) then grbp<="010";
	end if;
	if (ll=267 and cc>=29 and cc<42) then grbp<="010";
	end if;
	if (cc=46 and ll=267) then grbp<="010";
	end if;
	if (cc=66 and ll=267) then grbp<="010";
	end if;
	if (cc=81 and ll=267) then grbp<="010";
	end if;
	if (cc=106 and ll=267) then grbp<="010";
	end if;
	if (ll=267 and cc>=106 and cc<132) then grbp<="010";
	end if;
	if (ll=267 and cc>=136 and cc<153) then grbp<="010";
	end if;
	if (ll=267 and cc>=157 and cc<167) then grbp<="010";
	end if;
	if (cc=184 and ll=267) then grbp<="010";
	end if;
	if (ll=267 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=267 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (ll=267 and cc>=202 and cc<204) then grbp<="010";
	end if;
	if (ll=267 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=267 and cc>=214 and cc<224) then grbp<="010";
	end if;
	if (ll=268 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=268 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=268 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=55 and ll=268) then grbp<="010";
	end if;
	if (cc=79 and ll=268) then grbp<="010";
	end if;
	if (cc=96 and ll=268) then grbp<="010";
	end if;
	if (cc=106 and ll=268) then grbp<="010";
	end if;
	if (ll=268 and cc>=106 and cc<132) then grbp<="010";
	end if;
	if (ll=268 and cc>=136 and cc<145) then grbp<="010";
	end if;
	if (ll=268 and cc>=146 and cc<153) then grbp<="010";
	end if;
	if (ll=268 and cc>=157 and cc<167) then grbp<="010";
	end if;
	if (cc=176 and ll=268) then grbp<="010";
	end if;
	if (cc=184 and ll=268) then grbp<="010";
	end if;
	if (cc=186 and ll=268) then grbp<="010";
	end if;
	if (cc=190 and ll=268) then grbp<="010";
	end if;
	if (cc=192 and ll=268) then grbp<="010";
	end if;
	if (ll=268 and cc>=192 and cc<195) then grbp<="010";
	end if;
	if (ll=268 and cc>=205 and cc<207) then grbp<="010";
	end if;
	if (ll=268 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (cc=215 and ll=268) then grbp<="010";
	end if;
	if (cc=217 and ll=268) then grbp<="010";
	end if;
	if (ll=268 and cc>=217 and cc<224) then grbp<="010";
	end if;
	if (ll=269 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=269 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=269 and cc>=29 and cc<43) then grbp<="010";
	end if;
	if (cc=46 and ll=269) then grbp<="010";
	end if;
	if (ll=269 and cc>=46 and cc<48) then grbp<="010";
	end if;
	if (cc=70 and ll=269) then grbp<="010";
	end if;
	if (cc=79 and ll=269) then grbp<="010";
	end if;
	if (cc=106 and ll=269) then grbp<="010";
	end if;
	if (ll=269 and cc>=106 and cc<131) then grbp<="010";
	end if;
	if (ll=269 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (ll=269 and cc>=136 and cc<154) then grbp<="010";
	end if;
	if (ll=269 and cc>=158 and cc<166) then grbp<="010";
	end if;
	if (cc=176 and ll=269) then grbp<="010";
	end if;
	if (cc=182 and ll=269) then grbp<="010";
	end if;
	if (cc=184 and ll=269) then grbp<="010";
	end if;
	if (cc=186 and ll=269) then grbp<="010";
	end if;
	if (cc=190 and ll=269) then grbp<="010";
	end if;
	if (ll=269 and cc>=190 and cc<195) then grbp<="010";
	end if;
	if (cc=213 and ll=269) then grbp<="010";
	end if;
	if (ll=269 and cc>=213 and cc<224) then grbp<="010";
	end if;
	if (ll=270 and cc>=0 and cc<11) then grbp<="010";
	end if;
	if (ll=270 and cc>=12 and cc<17) then grbp<="010";
	end if;
	if (ll=270 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=48 and ll=270) then grbp<="010";
	end if;
	if (ll=270 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (cc=72 and ll=270) then grbp<="010";
	end if;
	if (cc=80 and ll=270) then grbp<="010";
	end if;
	if (cc=88 and ll=270) then grbp<="010";
	end if;
	if (ll=270 and cc>=88 and cc<90) then grbp<="010";
	end if;
	if (cc=105 and ll=270) then grbp<="010";
	end if;
	if (ll=270 and cc>=105 and cc<132) then grbp<="010";
	end if;
	if (ll=270 and cc>=136 and cc<154) then grbp<="010";
	end if;
	if (ll=270 and cc>=158 and cc<166) then grbp<="010";
	end if;
	if (cc=176 and ll=270) then grbp<="010";
	end if;
	if (cc=182 and ll=270) then grbp<="010";
	end if;
	if (cc=184 and ll=270) then grbp<="010";
	end if;
	if (cc=186 and ll=270) then grbp<="010";
	end if;
	if (cc=189 and ll=270) then grbp<="010";
	end if;
	if (ll=270 and cc>=189 and cc<195) then grbp<="010";
	end if;
	if (ll=270 and cc>=208 and cc<210) then grbp<="010";
	end if;
	if (ll=270 and cc>=211 and cc<224) then grbp<="010";
	end if;
	if (ll=271 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=271 and cc>=29 and cc<45) then grbp<="010";
	end if;
	if (cc=48 and ll=271) then grbp<="010";
	end if;
	if (cc=72 and ll=271) then grbp<="010";
	end if;
	if (ll=271 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=271 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=271 and cc>=105 and cc<133) then grbp<="010";
	end if;
	if (ll=271 and cc>=136 and cc<153) then grbp<="010";
	end if;
	if (ll=271 and cc>=158 and cc<166) then grbp<="010";
	end if;
	if (cc=176 and ll=271) then grbp<="010";
	end if;
	if (cc=182 and ll=271) then grbp<="010";
	end if;
	if (cc=185 and ll=271) then grbp<="010";
	end if;
	if (ll=271 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=271 and cc>=189 and cc<194) then grbp<="010";
	end if;
	if (cc=211 and ll=271) then grbp<="010";
	end if;
	if (ll=271 and cc>=211 and cc<216) then grbp<="010";
	end if;
	if (ll=271 and cc>=217 and cc<223) then grbp<="010";
	end if;
	if (ll=272 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=272 and cc>=29 and cc<44) then grbp<="010";
	end if;
	if (cc=73 and ll=272) then grbp<="010";
	end if;
	if (cc=84 and ll=272) then grbp<="010";
	end if;
	if (ll=272 and cc>=84 and cc<92) then grbp<="010";
	end if;
	if (cc=105 and ll=272) then grbp<="010";
	end if;
	if (ll=272 and cc>=105 and cc<133) then grbp<="010";
	end if;
	if (cc=137 and ll=272) then grbp<="010";
	end if;
	if (ll=272 and cc>=137 and cc<151) then grbp<="010";
	end if;
	if (ll=272 and cc>=158 and cc<166) then grbp<="010";
	end if;
	if (cc=176 and ll=272) then grbp<="010";
	end if;
	if (cc=182 and ll=272) then grbp<="010";
	end if;
	if (cc=185 and ll=272) then grbp<="010";
	end if;
	if (ll=272 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=272 and cc>=189 and cc<194) then grbp<="010";
	end if;
	if (cc=210 and ll=272) then grbp<="010";
	end if;
	if (cc=212 and ll=272) then grbp<="010";
	end if;
	if (cc=214 and ll=272) then grbp<="010";
	end if;
	if (ll=272 and cc>=214 and cc<223) then grbp<="010";
	end if;
	if (ll=273 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=273 and cc>=29 and cc<43) then grbp<="010";
	end if;
	if (cc=63 and ll=273) then grbp<="010";
	end if;
	if (cc=73 and ll=273) then grbp<="010";
	end if;
	if (ll=273 and cc>=73 and cc<75) then grbp<="010";
	end if;
	if (ll=273 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (ll=273 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=273 and cc>=105 and cc<132) then grbp<="010";
	end if;
	if (ll=273 and cc>=133 and cc<135) then grbp<="010";
	end if;
	if (ll=273 and cc>=138 and cc<150) then grbp<="010";
	end if;
	if (ll=273 and cc>=157 and cc<165) then grbp<="010";
	end if;
	if (cc=176 and ll=273) then grbp<="010";
	end if;
	if (cc=182 and ll=273) then grbp<="010";
	end if;
	if (cc=185 and ll=273) then grbp<="010";
	end if;
	if (ll=273 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=273 and cc>=189 and cc<194) then grbp<="010";
	end if;
	if (ll=273 and cc>=208 and cc<210) then grbp<="010";
	end if;
	if (ll=273 and cc>=211 and cc<213) then grbp<="010";
	end if;
	if (ll=273 and cc>=214 and cc<223) then grbp<="010";
	end if;
	if (ll=274 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=274 and cc>=29 and cc<43) then grbp<="010";
	end if;
	if (cc=52 and ll=274) then grbp<="010";
	end if;
	if (cc=67 and ll=274) then grbp<="010";
	end if;
	if (cc=72 and ll=274) then grbp<="010";
	end if;
	if (cc=74 and ll=274) then grbp<="010";
	end if;
	if (cc=78 and ll=274) then grbp<="010";
	end if;
	if (cc=82 and ll=274) then grbp<="010";
	end if;
	if (ll=274 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=274 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=274 and cc>=105 and cc<134) then grbp<="010";
	end if;
	if (ll=274 and cc>=136 and cc<150) then grbp<="010";
	end if;
	if (ll=274 and cc>=157 and cc<165) then grbp<="010";
	end if;
	if (cc=176 and ll=274) then grbp<="010";
	end if;
	if (cc=182 and ll=274) then grbp<="010";
	end if;
	if (cc=185 and ll=274) then grbp<="010";
	end if;
	if (ll=274 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=274 and cc>=189 and cc<194) then grbp<="010";
	end if;
	if (cc=210 and ll=274) then grbp<="010";
	end if;
	if (ll=274 and cc>=210 and cc<223) then grbp<="010";
	end if;
	if (ll=275 and cc>=0 and cc<17) then grbp<="010";
	end if;
	if (ll=275 and cc>=29 and cc<42) then grbp<="010";
	end if;
	if (ll=275 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=275 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (ll=275 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=105 and ll=275) then grbp<="010";
	end if;
	if (ll=275 and cc>=105 and cc<133) then grbp<="010";
	end if;
	if (ll=275 and cc>=135 and cc<138) then grbp<="010";
	end if;
	if (ll=275 and cc>=139 and cc<147) then grbp<="010";
	end if;
	if (cc=157 and ll=275) then grbp<="010";
	end if;
	if (ll=275 and cc>=157 and cc<165) then grbp<="010";
	end if;
	if (ll=275 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=182 and ll=275) then grbp<="010";
	end if;
	if (cc=185 and ll=275) then grbp<="010";
	end if;
	if (ll=275 and cc>=185 and cc<188) then grbp<="010";
	end if;
	if (ll=275 and cc>=189 and cc<194) then grbp<="010";
	end if;
	if (cc=206 and ll=275) then grbp<="010";
	end if;
	if (ll=275 and cc>=206 and cc<208) then grbp<="010";
	end if;
	if (ll=275 and cc>=211 and cc<223) then grbp<="010";
	end if;
	if (ll=276 and cc>=0 and cc<16) then grbp<="010";
	end if;
	if (ll=276 and cc>=29 and cc<42) then grbp<="010";
	end if;
	if (cc=51 and ll=276) then grbp<="010";
	end if;
	if (cc=72 and ll=276) then grbp<="010";
	end if;
	if (ll=276 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=276 and cc>=80 and cc<84) then grbp<="010";
	end if;
	if (ll=276 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (ll=276 and cc>=105 and cc<133) then grbp<="010";
	end if;
	if (cc=137 and ll=276) then grbp<="010";
	end if;
	if (ll=276 and cc>=137 and cc<147) then grbp<="010";
	end if;
	if (cc=157 and ll=276) then grbp<="010";
	end if;
	if (ll=276 and cc>=157 and cc<164) then grbp<="010";
	end if;
	if (ll=276 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=182 and ll=276) then grbp<="010";
	end if;
	if (cc=185 and ll=276) then grbp<="010";
	end if;
	if (ll=276 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (ll=276 and cc>=205 and cc<208) then grbp<="010";
	end if;
	if (cc=211 and ll=276) then grbp<="010";
	end if;
	if (ll=276 and cc>=211 and cc<214) then grbp<="010";
	end if;
	if (ll=276 and cc>=215 and cc<223) then grbp<="010";
	end if;
	if (ll=277 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=277 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=277 and cc>=29 and cc<41) then grbp<="010";
	end if;
	if (cc=46 and ll=277) then grbp<="010";
	end if;
	if (cc=72 and ll=277) then grbp<="010";
	end if;
	if (ll=277 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (cc=82 and ll=277) then grbp<="010";
	end if;
	if (cc=87 and ll=277) then grbp<="010";
	end if;
	if (ll=277 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (cc=106 and ll=277) then grbp<="010";
	end if;
	if (ll=277 and cc>=106 and cc<146) then grbp<="010";
	end if;
	if (ll=277 and cc>=157 and cc<164) then grbp<="010";
	end if;
	if (ll=277 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=182 and ll=277) then grbp<="010";
	end if;
	if (cc=185 and ll=277) then grbp<="010";
	end if;
	if (ll=277 and cc>=185 and cc<194) then grbp<="010";
	end if;
	if (cc=209 and ll=277) then grbp<="010";
	end if;
	if (ll=277 and cc>=209 and cc<213) then grbp<="010";
	end if;
	if (ll=277 and cc>=215 and cc<223) then grbp<="010";
	end if;
	if (ll=278 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=278 and cc>=11 and cc<16) then grbp<="010";
	end if;
	if (ll=278 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (ll=278 and cc>=42 and cc<44) then grbp<="010";
	end if;
	if (cc=68 and ll=278) then grbp<="010";
	end if;
	if (cc=70 and ll=278) then grbp<="010";
	end if;
	if (ll=278 and cc>=70 and cc<74) then grbp<="010";
	end if;
	if (ll=278 and cc>=86 and cc<90) then grbp<="010";
	end if;
	if (ll=278 and cc>=105 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=278) then grbp<="010";
	end if;
	if (ll=278 and cc>=137 and cc<146) then grbp<="010";
	end if;
	if (ll=278 and cc>=157 and cc<164) then grbp<="010";
	end if;
	if (cc=173 and ll=278) then grbp<="010";
	end if;
	if (ll=278 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=185 and ll=278) then grbp<="010";
	end if;
	if (ll=278 and cc>=185 and cc<190) then grbp<="010";
	end if;
	if (ll=278 and cc>=191 and cc<193) then grbp<="010";
	end if;
	if (cc=209 and ll=278) then grbp<="010";
	end if;
	if (ll=278 and cc>=209 and cc<212) then grbp<="010";
	end if;
	if (ll=278 and cc>=213 and cc<223) then grbp<="010";
	end if;
	if (ll=279 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=279 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=279 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (ll=279 and cc>=41 and cc<44) then grbp<="010";
	end if;
	if (ll=279 and cc>=70 and cc<74) then grbp<="010";
	end if;
	if (cc=86 and ll=279) then grbp<="010";
	end if;
	if (ll=279 and cc>=86 and cc<90) then grbp<="010";
	end if;
	if (cc=106 and ll=279) then grbp<="010";
	end if;
	if (ll=279 and cc>=106 and cc<136) then grbp<="010";
	end if;
	if (ll=279 and cc>=137 and cc<146) then grbp<="010";
	end if;
	if (ll=279 and cc>=157 and cc<163) then grbp<="010";
	end if;
	if (ll=279 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=185 and ll=279) then grbp<="010";
	end if;
	if (ll=279 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (cc=205 and ll=279) then grbp<="010";
	end if;
	if (cc=207 and ll=279) then grbp<="010";
	end if;
	if (ll=279 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=279 and cc>=210 and cc<215) then grbp<="010";
	end if;
	if (ll=279 and cc>=216 and cc<223) then grbp<="010";
	end if;
	if (ll=280 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=280 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=280 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (cc=70 and ll=280) then grbp<="010";
	end if;
	if (ll=280 and cc>=70 and cc<73) then grbp<="010";
	end if;
	if (ll=280 and cc>=86 and cc<90) then grbp<="010";
	end if;
	if (ll=280 and cc>=106 and cc<136) then grbp<="010";
	end if;
	if (ll=280 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=280 and cc>=157 and cc<163) then grbp<="010";
	end if;
	if (ll=280 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=183 and ll=280) then grbp<="010";
	end if;
	if (cc=185 and ll=280) then grbp<="010";
	end if;
	if (ll=280 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (cc=208 and ll=280) then grbp<="010";
	end if;
	if (ll=280 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=280 and cc>=214 and cc<222) then grbp<="010";
	end if;
	if (ll=281 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=281 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=281 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (ll=281 and cc>=40 and cc<43) then grbp<="010";
	end if;
	if (cc=70 and ll=281) then grbp<="010";
	end if;
	if (ll=281 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (ll=281 and cc>=77 and cc<81) then grbp<="010";
	end if;
	if (ll=281 and cc>=85 and cc<89) then grbp<="010";
	end if;
	if (cc=106 and ll=281) then grbp<="010";
	end if;
	if (ll=281 and cc>=106 and cc<145) then grbp<="010";
	end if;
	if (ll=281 and cc>=157 and cc<163) then grbp<="010";
	end if;
	if (ll=281 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=183 and ll=281) then grbp<="010";
	end if;
	if (cc=185 and ll=281) then grbp<="010";
	end if;
	if (ll=281 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (cc=205 and ll=281) then grbp<="010";
	end if;
	if (cc=208 and ll=281) then grbp<="010";
	end if;
	if (ll=281 and cc>=208 and cc<222) then grbp<="010";
	end if;
	if (ll=282 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=282 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=282 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (ll=282 and cc>=40 and cc<43) then grbp<="010";
	end if;
	if (cc=69 and ll=282) then grbp<="010";
	end if;
	if (ll=282 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=282 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=282 and cc>=85 and cc<89) then grbp<="010";
	end if;
	if (ll=282 and cc>=106 and cc<145) then grbp<="010";
	end if;
	if (ll=282 and cc>=156 and cc<163) then grbp<="010";
	end if;
	if (ll=282 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=183 and ll=282) then grbp<="010";
	end if;
	if (cc=185 and ll=282) then grbp<="010";
	end if;
	if (ll=282 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (ll=282 and cc>=201 and cc<203) then grbp<="010";
	end if;
	if (cc=208 and ll=282) then grbp<="010";
	end if;
	if (ll=282 and cc>=208 and cc<211) then grbp<="010";
	end if;
	if (cc=214 and ll=282) then grbp<="010";
	end if;
	if (ll=282 and cc>=214 and cc<222) then grbp<="010";
	end if;
	if (ll=283 and cc>=0 and cc<9) then grbp<="010";
	end if;
	if (ll=283 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=283 and cc>=29 and cc<38) then grbp<="010";
	end if;
	if (ll=283 and cc>=39 and cc<43) then grbp<="010";
	end if;
	if (cc=57 and ll=283) then grbp<="010";
	end if;
	if (cc=71 and ll=283) then grbp<="010";
	end if;
	if (cc=75 and ll=283) then grbp<="010";
	end if;
	if (ll=283 and cc>=75 and cc<80) then grbp<="010";
	end if;
	if (ll=283 and cc>=84 and cc<88) then grbp<="010";
	end if;
	if (ll=283 and cc>=106 and cc<144) then grbp<="010";
	end if;
	if (ll=283 and cc>=156 and cc<162) then grbp<="010";
	end if;
	if (ll=283 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (cc=185 and ll=283) then grbp<="010";
	end if;
	if (ll=283 and cc>=185 and cc<193) then grbp<="010";
	end if;
	if (cc=207 and ll=283) then grbp<="010";
	end if;
	if (ll=283 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=283 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=283 and cc>=214 and cc<222) then grbp<="010";
	end if;
	if (ll=284 and cc>=0 and cc<8) then grbp<="010";
	end if;
	if (ll=284 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=284 and cc>=29 and cc<38) then grbp<="010";
	end if;
	if (ll=284 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=284 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=71 and ll=284) then grbp<="010";
	end if;
	if (cc=75 and ll=284) then grbp<="010";
	end if;
	if (ll=284 and cc>=75 and cc<80) then grbp<="010";
	end if;
	if (ll=284 and cc>=84 and cc<88) then grbp<="010";
	end if;
	if (cc=106 and ll=284) then grbp<="010";
	end if;
	if (ll=284 and cc>=106 and cc<145) then grbp<="010";
	end if;
	if (ll=284 and cc>=156 and cc<162) then grbp<="010";
	end if;
	if (ll=284 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (cc=185 and ll=284) then grbp<="010";
	end if;
	if (ll=284 and cc>=185 and cc<192) then grbp<="010";
	end if;
	if (cc=205 and ll=284) then grbp<="010";
	end if;
	if (cc=207 and ll=284) then grbp<="010";
	end if;
	if (ll=284 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=284 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (ll=284 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (cc=2 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=2 and cc<9) then grbp<="010";
	end if;
	if (ll=285 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=285 and cc>=29 and cc<37) then grbp<="010";
	end if;
	if (ll=285 and cc>=38 and cc<43) then grbp<="010";
	end if;
	if (cc=46 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=46 and cc<48) then grbp<="010";
	end if;
	if (cc=78 and ll=285) then grbp<="010";
	end if;
	if (cc=84 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=84 and cc<88) then grbp<="010";
	end if;
	if (cc=101 and ll=285) then grbp<="010";
	end if;
	if (cc=106 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=106 and cc<143) then grbp<="010";
	end if;
	if (ll=285 and cc>=156 and cc<162) then grbp<="010";
	end if;
	if (ll=285 and cc>=172 and cc<176) then grbp<="010";
	end if;
	if (cc=185 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=185 and cc<192) then grbp<="010";
	end if;
	if (ll=285 and cc>=202 and cc<204) then grbp<="010";
	end if;
	if (cc=207 and ll=285) then grbp<="010";
	end if;
	if (ll=285 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=285 and cc>=210 and cc<222) then grbp<="010";
	end if;
	if (cc=4 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=4 and cc<9) then grbp<="010";
	end if;
	if (ll=286 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=286 and cc>=29 and cc<37) then grbp<="010";
	end if;
	if (ll=286 and cc>=38 and cc<43) then grbp<="010";
	end if;
	if (cc=63 and ll=286) then grbp<="010";
	end if;
	if (cc=74 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=286 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (cc=93 and ll=286) then grbp<="010";
	end if;
	if (cc=101 and ll=286) then grbp<="010";
	end if;
	if (cc=106 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=106 and cc<142) then grbp<="010";
	end if;
	if (cc=156 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=156 and cc<162) then grbp<="010";
	end if;
	if (ll=286 and cc>=173 and cc<178) then grbp<="010";
	end if;
	if (cc=185 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=185 and cc<192) then grbp<="010";
	end if;
	if (cc=208 and ll=286) then grbp<="010";
	end if;
	if (ll=286 and cc>=208 and cc<222) then grbp<="010";
	end if;
	if (cc=4 and ll=287) then grbp<="010";
	end if;
	if (ll=287 and cc>=4 and cc<9) then grbp<="010";
	end if;
	if (ll=287 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=287 and cc>=29 and cc<43) then grbp<="010";
	end if;
	if (cc=68 and ll=287) then grbp<="010";
	end if;
	if (cc=74 and ll=287) then grbp<="010";
	end if;
	if (ll=287 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=287 and cc>=83 and cc<87) then grbp<="010";
	end if;
	if (cc=106 and ll=287) then grbp<="010";
	end if;
	if (ll=287 and cc>=106 and cc<149) then grbp<="010";
	end if;
	if (ll=287 and cc>=153 and cc<161) then grbp<="010";
	end if;
	if (ll=287 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=185 and ll=287) then grbp<="010";
	end if;
	if (ll=287 and cc>=185 and cc<192) then grbp<="010";
	end if;
	if (ll=287 and cc>=201 and cc<204) then grbp<="010";
	end if;
	if (ll=287 and cc>=206 and cc<208) then grbp<="010";
	end if;
	if (ll=287 and cc>=210 and cc<222) then grbp<="010";
	end if;
	if (cc=5 and ll=288) then grbp<="010";
	end if;
	if (ll=288 and cc>=5 and cc<9) then grbp<="010";
	end if;
	if (ll=288 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=288 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=288 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=46 and ll=288) then grbp<="010";
	end if;
	if (cc=58 and ll=288) then grbp<="010";
	end if;
	if (cc=73 and ll=288) then grbp<="010";
	end if;
	if (ll=288 and cc>=73 and cc<76) then grbp<="010";
	end if;
	if (ll=288 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (cc=100 and ll=288) then grbp<="010";
	end if;
	if (cc=106 and ll=288) then grbp<="010";
	end if;
	if (ll=288 and cc>=106 and cc<161) then grbp<="010";
	end if;
	if (ll=288 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=185 and ll=288) then grbp<="010";
	end if;
	if (ll=288 and cc>=185 and cc<192) then grbp<="010";
	end if;
	if (ll=288 and cc>=201 and cc<204) then grbp<="010";
	end if;
	if (cc=209 and ll=288) then grbp<="010";
	end if;
	if (ll=288 and cc>=209 and cc<213) then grbp<="010";
	end if;
	if (ll=288 and cc>=214 and cc<222) then grbp<="010";
	end if;
	if (ll=289 and cc>=6 and cc<8) then grbp<="010";
	end if;
	if (ll=289 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=289 and cc>=29 and cc<41) then grbp<="010";
	end if;
	if (cc=47 and ll=289) then grbp<="010";
	end if;
	if (cc=58 and ll=289) then grbp<="010";
	end if;
	if (ll=289 and cc>=58 and cc<60) then grbp<="010";
	end if;
	if (ll=289 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (cc=102 and ll=289) then grbp<="010";
	end if;
	if (cc=106 and ll=289) then grbp<="010";
	end if;
	if (ll=289 and cc>=106 and cc<161) then grbp<="010";
	end if;
	if (ll=289 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=185 and ll=289) then grbp<="010";
	end if;
	if (cc=187 and ll=289) then grbp<="010";
	end if;
	if (ll=289 and cc>=187 and cc<192) then grbp<="010";
	end if;
	if (cc=207 and ll=289) then grbp<="010";
	end if;
	if (cc=209 and ll=289) then grbp<="010";
	end if;
	if (ll=289 and cc>=209 and cc<222) then grbp<="010";
	end if;
	if (cc=10 and ll=290) then grbp<="010";
	end if;
	if (ll=290 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=290 and cc>=29 and cc<35) then grbp<="010";
	end if;
	if (ll=290 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (cc=81 and ll=290) then grbp<="010";
	end if;
	if (ll=290 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (cc=102 and ll=290) then grbp<="010";
	end if;
	if (cc=106 and ll=290) then grbp<="010";
	end if;
	if (ll=290 and cc>=106 and cc<160) then grbp<="010";
	end if;
	if (ll=290 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=187 and ll=290) then grbp<="010";
	end if;
	if (ll=290 and cc>=187 and cc<192) then grbp<="010";
	end if;
	if (cc=207 and ll=290) then grbp<="010";
	end if;
	if (ll=290 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=290 and cc>=211 and cc<222) then grbp<="010";
	end if;
	if (ll=291 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=291 and cc>=29 and cc<35) then grbp<="010";
	end if;
	if (ll=291 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (cc=72 and ll=291) then grbp<="010";
	end if;
	if (cc=74 and ll=291) then grbp<="010";
	end if;
	if (ll=291 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=291 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (cc=102 and ll=291) then grbp<="010";
	end if;
	if (cc=106 and ll=291) then grbp<="010";
	end if;
	if (ll=291 and cc>=106 and cc<160) then grbp<="010";
	end if;
	if (ll=291 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=183 and ll=291) then grbp<="010";
	end if;
	if (cc=186 and ll=291) then grbp<="010";
	end if;
	if (ll=291 and cc>=186 and cc<192) then grbp<="010";
	end if;
	if (cc=207 and ll=291) then grbp<="010";
	end if;
	if (cc=210 and ll=291) then grbp<="010";
	end if;
	if (ll=291 and cc>=210 and cc<222) then grbp<="010";
	end if;
	if (ll=292 and cc>=9 and cc<16) then grbp<="010";
	end if;
	if (ll=292 and cc>=29 and cc<34) then grbp<="010";
	end if;
	if (ll=292 and cc>=35 and cc<39) then grbp<="010";
	end if;
	if (cc=72 and ll=292) then grbp<="010";
	end if;
	if (ll=292 and cc>=72 and cc<76) then grbp<="010";
	end if;
	if (ll=292 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (cc=106 and ll=292) then grbp<="010";
	end if;
	if (ll=292 and cc>=106 and cc<160) then grbp<="010";
	end if;
	if (ll=292 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (cc=183 and ll=292) then grbp<="010";
	end if;
	if (cc=186 and ll=292) then grbp<="010";
	end if;
	if (ll=292 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (ll=292 and cc>=189 and cc<192) then grbp<="010";
	end if;
	if (cc=206 and ll=292) then grbp<="010";
	end if;
	if (cc=210 and ll=292) then grbp<="010";
	end if;
	if (ll=292 and cc>=210 and cc<222) then grbp<="010";
	end if;
	if (cc=8 and ll=293) then grbp<="010";
	end if;
	if (ll=293 and cc>=8 and cc<16) then grbp<="010";
	end if;
	if (ll=293 and cc>=29 and cc<34) then grbp<="010";
	end if;
	if (ll=293 and cc>=35 and cc<39) then grbp<="010";
	end if;
	if (ll=293 and cc>=41 and cc<43) then grbp<="010";
	end if;
	if (ll=293 and cc>=72 and cc<77) then grbp<="010";
	end if;
	if (ll=293 and cc>=80 and cc<84) then grbp<="010";
	end if;
	if (cc=106 and ll=293) then grbp<="010";
	end if;
	if (ll=293 and cc>=106 and cc<148) then grbp<="010";
	end if;
	if (ll=293 and cc>=152 and cc<159) then grbp<="010";
	end if;
	if (ll=293 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=293) then grbp<="010";
	end if;
	if (cc=186 and ll=293) then grbp<="010";
	end if;
	if (ll=293 and cc>=186 and cc<191) then grbp<="010";
	end if;
	if (cc=206 and ll=293) then grbp<="010";
	end if;
	if (cc=210 and ll=293) then grbp<="010";
	end if;
	if (cc=212 and ll=293) then grbp<="010";
	end if;
	if (ll=293 and cc>=212 and cc<222) then grbp<="010";
	end if;
	if (ll=294 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=294 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=294 and cc>=34 and cc<39) then grbp<="010";
	end if;
	if (ll=294 and cc>=40 and cc<43) then grbp<="010";
	end if;
	if (cc=65 and ll=294) then grbp<="010";
	end if;
	if (ll=294 and cc>=65 and cc<67) then grbp<="010";
	end if;
	if (ll=294 and cc>=73 and cc<77) then grbp<="010";
	end if;
	if (ll=294 and cc>=80 and cc<83) then grbp<="010";
	end if;
	if (cc=102 and ll=294) then grbp<="010";
	end if;
	if (cc=106 and ll=294) then grbp<="010";
	end if;
	if (cc=108 and ll=294) then grbp<="010";
	end if;
	if (ll=294 and cc>=108 and cc<143) then grbp<="010";
	end if;
	if (ll=294 and cc>=152 and cc<159) then grbp<="010";
	end if;
	if (ll=294 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=294) then grbp<="010";
	end if;
	if (cc=186 and ll=294) then grbp<="010";
	end if;
	if (ll=294 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (ll=294 and cc>=189 and cc<191) then grbp<="010";
	end if;
	if (cc=205 and ll=294) then grbp<="010";
	end if;
	if (ll=294 and cc>=205 and cc<208) then grbp<="010";
	end if;
	if (cc=211 and ll=294) then grbp<="010";
	end if;
	if (ll=294 and cc>=211 and cc<222) then grbp<="010";
	end if;
	if (ll=295 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=295 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (ll=295 and cc>=34 and cc<39) then grbp<="010";
	end if;
	if (ll=295 and cc>=40 and cc<43) then grbp<="010";
	end if;
	if (ll=295 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=295 and cc>=73 and cc<77) then grbp<="010";
	end if;
	if (ll=295 and cc>=79 and cc<83) then grbp<="010";
	end if;
	if (cc=108 and ll=295) then grbp<="010";
	end if;
	if (ll=295 and cc>=108 and cc<142) then grbp<="010";
	end if;
	if (ll=295 and cc>=152 and cc<159) then grbp<="010";
	end if;
	if (ll=295 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (cc=186 and ll=295) then grbp<="010";
	end if;
	if (ll=295 and cc>=186 and cc<191) then grbp<="010";
	end if;
	if (ll=295 and cc>=209 and cc<212) then grbp<="010";
	end if;
	if (ll=295 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=296 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=296 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (ll=296 and cc>=33 and cc<38) then grbp<="010";
	end if;
	if (ll=296 and cc>=39 and cc<43) then grbp<="010";
	end if;
	if (ll=296 and cc>=73 and cc<77) then grbp<="010";
	end if;
	if (ll=296 and cc>=79 and cc<82) then grbp<="010";
	end if;
	if (cc=106 and ll=296) then grbp<="010";
	end if;
	if (cc=108 and ll=296) then grbp<="010";
	end if;
	if (ll=296 and cc>=108 and cc<142) then grbp<="010";
	end if;
	if (ll=296 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (ll=296 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (cc=186 and ll=296) then grbp<="010";
	end if;
	if (ll=296 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (cc=207 and ll=296) then grbp<="010";
	end if;
	if (cc=209 and ll=296) then grbp<="010";
	end if;
	if (ll=296 and cc>=209 and cc<212) then grbp<="010";
	end if;
	if (ll=296 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=297 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=297 and cc>=33 and cc<38) then grbp<="010";
	end if;
	if (ll=297 and cc>=39 and cc<43) then grbp<="010";
	end if;
	if (cc=74 and ll=297) then grbp<="010";
	end if;
	if (ll=297 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=297 and cc>=78 and cc<81) then grbp<="010";
	end if;
	if (cc=106 and ll=297) then grbp<="010";
	end if;
	if (cc=108 and ll=297) then grbp<="010";
	end if;
	if (ll=297 and cc>=108 and cc<144) then grbp<="010";
	end if;
	if (ll=297 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (ll=297 and cc>=172 and cc<176) then grbp<="010";
	end if;
	if (cc=184 and ll=297) then grbp<="010";
	end if;
	if (cc=186 and ll=297) then grbp<="010";
	end if;
	if (ll=297 and cc>=186 and cc<188) then grbp<="010";
	end if;
	if (cc=209 and ll=297) then grbp<="010";
	end if;
	if (ll=297 and cc>=209 and cc<212) then grbp<="010";
	end if;
	if (ll=297 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=298 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=298 and cc>=32 and cc<37) then grbp<="010";
	end if;
	if (ll=298 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=298 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=298 and cc>=78 and cc<81) then grbp<="010";
	end if;
	if (cc=108 and ll=298) then grbp<="010";
	end if;
	if (ll=298 and cc>=108 and cc<144) then grbp<="010";
	end if;
	if (cc=151 and ll=298) then grbp<="010";
	end if;
	if (ll=298 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (ll=298 and cc>=172 and cc<176) then grbp<="010";
	end if;
	if (cc=184 and ll=298) then grbp<="010";
	end if;
	if (cc=186 and ll=298) then grbp<="010";
	end if;
	if (cc=189 and ll=298) then grbp<="010";
	end if;
	if (ll=298 and cc>=189 and cc<192) then grbp<="010";
	end if;
	if (ll=298 and cc>=209 and cc<222) then grbp<="010";
	end if;
	if (ll=299 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=299 and cc>=31 and cc<37) then grbp<="010";
	end if;
	if (ll=299 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (ll=299 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=299 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (cc=108 and ll=299) then grbp<="010";
	end if;
	if (cc=110 and ll=299) then grbp<="010";
	end if;
	if (ll=299 and cc>=110 and cc<145) then grbp<="010";
	end if;
	if (ll=299 and cc>=147 and cc<158) then grbp<="010";
	end if;
	if (cc=174 and ll=299) then grbp<="010";
	end if;
	if (ll=299 and cc>=174 and cc<177) then grbp<="010";
	end if;
	if (cc=186 and ll=299) then grbp<="010";
	end if;
	if (cc=189 and ll=299) then grbp<="010";
	end if;
	if (cc=208 and ll=299) then grbp<="010";
	end if;
	if (ll=299 and cc>=208 and cc<211) then grbp<="010";
	end if;
	if (ll=299 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=300 and cc>=10 and cc<16) then grbp<="010";
	end if;
	if (ll=300 and cc>=30 and cc<37) then grbp<="010";
	end if;
	if (ll=300 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (cc=70 and ll=300) then grbp<="010";
	end if;
	if (cc=74 and ll=300) then grbp<="010";
	end if;
	if (ll=300 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (ll=300 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (cc=106 and ll=300) then grbp<="010";
	end if;
	if (cc=108 and ll=300) then grbp<="010";
	end if;
	if (cc=111 and ll=300) then grbp<="010";
	end if;
	if (ll=300 and cc>=111 and cc<157) then grbp<="010";
	end if;
	if (cc=174 and ll=300) then grbp<="010";
	end if;
	if (ll=300 and cc>=174 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=300) then grbp<="010";
	end if;
	if (cc=186 and ll=300) then grbp<="010";
	end if;
	if (cc=189 and ll=300) then grbp<="010";
	end if;
	if (cc=209 and ll=300) then grbp<="010";
	end if;
	if (ll=300 and cc>=209 and cc<222) then grbp<="010";
	end if;
	if (ll=301 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=301 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=301 and cc>=37 and cc<42) then grbp<="010";
	end if;
	if (ll=301 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (cc=108 and ll=301) then grbp<="010";
	end if;
	if (ll=301 and cc>=108 and cc<110) then grbp<="010";
	end if;
	if (ll=301 and cc>=111 and cc<157) then grbp<="010";
	end if;
	if (cc=174 and ll=301) then grbp<="010";
	end if;
	if (ll=301 and cc>=174 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=301) then grbp<="010";
	end if;
	if (cc=186 and ll=301) then grbp<="010";
	end if;
	if (cc=189 and ll=301) then grbp<="010";
	end if;
	if (cc=209 and ll=301) then grbp<="010";
	end if;
	if (ll=301 and cc>=209 and cc<222) then grbp<="010";
	end if;
	if (ll=302 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=302 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=302 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=71 and ll=302) then grbp<="010";
	end if;
	if (cc=75 and ll=302) then grbp<="010";
	end if;
	if (cc=81 and ll=302) then grbp<="010";
	end if;
	if (cc=108 and ll=302) then grbp<="010";
	end if;
	if (ll=302 and cc>=108 and cc<110) then grbp<="010";
	end if;
	if (ll=302 and cc>=111 and cc<157) then grbp<="010";
	end if;
	if (ll=302 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (ll=302 and cc>=179 and cc<181) then grbp<="010";
	end if;
	if (cc=186 and ll=302) then grbp<="010";
	end if;
	if (cc=189 and ll=302) then grbp<="010";
	end if;
	if (cc=210 and ll=302) then grbp<="010";
	end if;
	if (cc=212 and ll=302) then grbp<="010";
	end if;
	if (ll=302 and cc>=212 and cc<222) then grbp<="010";
	end if;
	if (ll=303 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=303 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=303 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=69 and ll=303) then grbp<="010";
	end if;
	if (cc=73 and ll=303) then grbp<="010";
	end if;
	if (cc=107 and ll=303) then grbp<="010";
	end if;
	if (ll=303 and cc>=107 and cc<110) then grbp<="010";
	end if;
	if (ll=303 and cc>=112 and cc<157) then grbp<="010";
	end if;
	if (ll=303 and cc>=171 and cc<177) then grbp<="010";
	end if;
	if (cc=184 and ll=303) then grbp<="010";
	end if;
	if (cc=186 and ll=303) then grbp<="010";
	end if;
	if (cc=189 and ll=303) then grbp<="010";
	end if;
	if (ll=303 and cc>=189 and cc<191) then grbp<="010";
	end if;
	if (ll=303 and cc>=209 and cc<212) then grbp<="010";
	end if;
	if (ll=303 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=304 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=304 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=304 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=50 and ll=304) then grbp<="010";
	end if;
	if (cc=70 and ll=304) then grbp<="010";
	end if;
	if (cc=73 and ll=304) then grbp<="010";
	end if;
	if (cc=77 and ll=304) then grbp<="010";
	end if;
	if (cc=80 and ll=304) then grbp<="010";
	end if;
	if (cc=109 and ll=304) then grbp<="010";
	end if;
	if (cc=112 and ll=304) then grbp<="010";
	end if;
	if (ll=304 and cc>=112 and cc<155) then grbp<="010";
	end if;
	if (cc=172 and ll=304) then grbp<="010";
	end if;
	if (ll=304 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (ll=304 and cc>=179 and cc<181) then grbp<="010";
	end if;
	if (cc=186 and ll=304) then grbp<="010";
	end if;
	if (cc=189 and ll=304) then grbp<="010";
	end if;
	if (cc=210 and ll=304) then grbp<="010";
	end if;
	if (ll=304 and cc>=210 and cc<222) then grbp<="010";
	end if;
	if (ll=305 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=305 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=305 and cc>=37 and cc<40) then grbp<="010";
	end if;
	if (cc=73 and ll=305) then grbp<="010";
	end if;
	if (cc=75 and ll=305) then grbp<="010";
	end if;
	if (cc=109 and ll=305) then grbp<="010";
	end if;
	if (cc=112 and ll=305) then grbp<="010";
	end if;
	if (ll=305 and cc>=112 and cc<155) then grbp<="010";
	end if;
	if (cc=172 and ll=305) then grbp<="010";
	end if;
	if (ll=305 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (ll=305 and cc>=179 and cc<181) then grbp<="010";
	end if;
	if (cc=189 and ll=305) then grbp<="010";
	end if;
	if (cc=212 and ll=305) then grbp<="010";
	end if;
	if (ll=305 and cc>=212 and cc<222) then grbp<="010";
	end if;
	if (ll=306 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=306 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=306 and cc>=37 and cc<40) then grbp<="010";
	end if;
	if (ll=306 and cc>=112 and cc<148) then grbp<="010";
	end if;
	if (ll=306 and cc>=149 and cc<155) then grbp<="010";
	end if;
	if (cc=172 and ll=306) then grbp<="010";
	end if;
	if (ll=306 and cc>=172 and cc<177) then grbp<="010";
	end if;
	if (ll=306 and cc>=179 and cc<181) then grbp<="010";
	end if;
	if (cc=188 and ll=306) then grbp<="010";
	end if;
	if (ll=306 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=306 and cc>=211 and cc<222) then grbp<="010";
	end if;
	if (ll=307 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=307 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=307 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=73 and ll=307) then grbp<="010";
	end if;
	if (cc=79 and ll=307) then grbp<="010";
	end if;
	if (cc=113 and ll=307) then grbp<="010";
	end if;
	if (ll=307 and cc>=113 and cc<142) then grbp<="010";
	end if;
	if (ll=307 and cc>=146 and cc<148) then grbp<="010";
	end if;
	if (ll=307 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (cc=172 and ll=307) then grbp<="010";
	end if;
	if (ll=307 and cc>=172 and cc<181) then grbp<="010";
	end if;
	if (cc=188 and ll=307) then grbp<="010";
	end if;
	if (ll=307 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (cc=213 and ll=307) then grbp<="010";
	end if;
	if (ll=307 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=308 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=308 and cc>=29 and cc<36) then grbp<="010";
	end if;
	if (ll=308 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (cc=70 and ll=308) then grbp<="010";
	end if;
	if (ll=308 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=113 and ll=308) then grbp<="010";
	end if;
	if (ll=308 and cc>=113 and cc<141) then grbp<="010";
	end if;
	if (cc=149 and ll=308) then grbp<="010";
	end if;
	if (ll=308 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=308 and cc>=172 and cc<181) then grbp<="010";
	end if;
	if (cc=188 and ll=308) then grbp<="010";
	end if;
	if (ll=308 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=308 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (ll=308 and cc>=213 and cc<222) then grbp<="010";
	end if;
	if (ll=309 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=309 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (ll=309 and cc>=42 and cc<44) then grbp<="010";
	end if;
	if (ll=309 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=78 and ll=309) then grbp<="010";
	end if;
	if (cc=113 and ll=309) then grbp<="010";
	end if;
	if (ll=309 and cc>=113 and cc<141) then grbp<="010";
	end if;
	if (cc=149 and ll=309) then grbp<="010";
	end if;
	if (ll=309 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=309 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=188 and ll=309) then grbp<="010";
	end if;
	if (cc=210 and ll=309) then grbp<="010";
	end if;
	if (cc=212 and ll=309) then grbp<="010";
	end if;
	if (ll=309 and cc>=212 and cc<222) then grbp<="010";
	end if;
	if (ll=310 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=310 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (ll=310 and cc>=42 and cc<44) then grbp<="010";
	end if;
	if (ll=310 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=113 and ll=310) then grbp<="010";
	end if;
	if (cc=116 and ll=310) then grbp<="010";
	end if;
	if (ll=310 and cc>=116 and cc<137) then grbp<="010";
	end if;
	if (ll=310 and cc>=138 and cc<140) then grbp<="010";
	end if;
	if (ll=310 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=310 and cc>=171 and cc<177) then grbp<="010";
	end if;
	if (ll=310 and cc>=178 and cc<180) then grbp<="010";
	end if;
	if (cc=188 and ll=310) then grbp<="010";
	end if;
	if (cc=210 and ll=310) then grbp<="010";
	end if;
	if (ll=310 and cc>=210 and cc<212) then grbp<="010";
	end if;
	if (ll=310 and cc>=213 and cc<221) then grbp<="010";
	end if;
	if (ll=311 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=311 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (cc=70 and ll=311) then grbp<="010";
	end if;
	if (ll=311 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=113 and ll=311) then grbp<="010";
	end if;
	if (cc=116 and ll=311) then grbp<="010";
	end if;
	if (ll=311 and cc>=116 and cc<136) then grbp<="010";
	end if;
	if (ll=311 and cc>=150 and cc<154) then grbp<="010";
	end if;
	if (ll=311 and cc>=171 and cc<177) then grbp<="010";
	end if;
	if (ll=311 and cc>=178 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=311) then grbp<="010";
	end if;
	if (cc=188 and ll=311) then grbp<="010";
	end if;
	if (ll=311 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=311 and cc>=211 and cc<221) then grbp<="010";
	end if;
	if (ll=312 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=312 and cc>=29 and cc<40) then grbp<="010";
	end if;
	if (cc=56 and ll=312) then grbp<="010";
	end if;
	if (cc=70 and ll=312) then grbp<="010";
	end if;
	if (ll=312 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=113 and ll=312) then grbp<="010";
	end if;
	if (cc=117 and ll=312) then grbp<="010";
	end if;
	if (ll=312 and cc>=117 and cc<136) then grbp<="010";
	end if;
	if (ll=312 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (cc=171 and ll=312) then grbp<="010";
	end if;
	if (ll=312 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=312) then grbp<="010";
	end if;
	if (cc=188 and ll=312) then grbp<="010";
	end if;
	if (cc=196 and ll=312) then grbp<="010";
	end if;
	if (cc=210 and ll=312) then grbp<="010";
	end if;
	if (ll=312 and cc>=210 and cc<221) then grbp<="010";
	end if;
	if (ll=313 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=313 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (cc=71 and ll=313) then grbp<="010";
	end if;
	if (cc=75 and ll=313) then grbp<="010";
	end if;
	if (ll=313 and cc>=75 and cc<78) then grbp<="010";
	end if;
	if (ll=313 and cc>=113 and cc<115) then grbp<="010";
	end if;
	if (ll=313 and cc>=118 and cc<135) then grbp<="010";
	end if;
	if (ll=313 and cc>=150 and cc<153) then grbp<="010";
	end if;
	if (ll=313 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=313) then grbp<="010";
	end if;
	if (cc=188 and ll=313) then grbp<="010";
	end if;
	if (cc=206 and ll=313) then grbp<="010";
	end if;
	if (cc=208 and ll=313) then grbp<="010";
	end if;
	if (cc=210 and ll=313) then grbp<="010";
	end if;
	if (ll=313 and cc>=210 and cc<221) then grbp<="010";
	end if;
	if (ll=314 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=314 and cc>=29 and cc<39) then grbp<="010";
	end if;
	if (cc=75 and ll=314) then grbp<="010";
	end if;
	if (cc=113 and ll=314) then grbp<="010";
	end if;
	if (ll=314 and cc>=113 and cc<115) then grbp<="010";
	end if;
	if (ll=314 and cc>=119 and cc<137) then grbp<="010";
	end if;
	if (ll=314 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=314 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=314) then grbp<="010";
	end if;
	if (cc=188 and ll=314) then grbp<="010";
	end if;
	if (cc=210 and ll=314) then grbp<="010";
	end if;
	if (ll=314 and cc>=210 and cc<221) then grbp<="010";
	end if;
	if (ll=315 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=315 and cc>=29 and cc<38) then grbp<="010";
	end if;
	if (ll=315 and cc>=73 and cc<76) then grbp<="010";
	end if;
	if (ll=315 and cc>=113 and cc<115) then grbp<="010";
	end if;
	if (ll=315 and cc>=119 and cc<138) then grbp<="010";
	end if;
	if (ll=315 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=315 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=315) then grbp<="010";
	end if;
	if (cc=188 and ll=315) then grbp<="010";
	end if;
	if (cc=196 and ll=315) then grbp<="010";
	end if;
	if (cc=208 and ll=315) then grbp<="010";
	end if;
	if (ll=315 and cc>=208 and cc<221) then grbp<="010";
	end if;
	if (ll=316 and cc>=9 and cc<17) then grbp<="010";
	end if;
	if (ll=316 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=316 and cc>=35 and cc<38) then grbp<="010";
	end if;
	if (cc=73 and ll=316) then grbp<="010";
	end if;
	if (ll=316 and cc>=73 and cc<76) then grbp<="010";
	end if;
	if (cc=120 and ll=316) then grbp<="010";
	end if;
	if (ll=316 and cc>=120 and cc<138) then grbp<="010";
	end if;
	if (ll=316 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=316 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=316) then grbp<="010";
	end if;
	if (cc=188 and ll=316) then grbp<="010";
	end if;
	if (cc=208 and ll=316) then grbp<="010";
	end if;
	if (cc=210 and ll=316) then grbp<="010";
	end if;
	if (ll=316 and cc>=210 and cc<221) then grbp<="010";
	end if;
	if (ll=316 and cc>=249 and cc<251) then grbp<="010";
	end if;
	if (cc=9 and ll=317) then grbp<="010";
	end if;
	if (ll=317 and cc>=9 and cc<18) then grbp<="010";
	end if;
	if (ll=317 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=317 and cc>=35 and cc<38) then grbp<="010";
	end if;
	if (ll=317 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=317 and cc>=75 and cc<77) then grbp<="010";
	end if;
	if (cc=115 and ll=317) then grbp<="010";
	end if;
	if (cc=121 and ll=317) then grbp<="010";
	end if;
	if (ll=317 and cc>=121 and cc<136) then grbp<="010";
	end if;
	if (cc=148 and ll=317) then grbp<="010";
	end if;
	if (ll=317 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=317 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=317) then grbp<="010";
	end if;
	if (cc=188 and ll=317) then grbp<="010";
	end if;
	if (ll=317 and cc>=188 and cc<191) then grbp<="010";
	end if;
	if (cc=204 and ll=317) then grbp<="010";
	end if;
	if (cc=207 and ll=317) then grbp<="010";
	end if;
	if (cc=209 and ll=317) then grbp<="010";
	end if;
	if (cc=211 and ll=317) then grbp<="010";
	end if;
	if (ll=317 and cc>=211 and cc<221) then grbp<="010";
	end if;
	if (ll=317 and cc>=247 and cc<250) then grbp<="010";
	end if;
	if (ll=318 and cc>=10 and cc<18) then grbp<="010";
	end if;
	if (ll=318 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=318 and cc>=35 and cc<38) then grbp<="010";
	end if;
	if (cc=58 and ll=318) then grbp<="010";
	end if;
	if (cc=76 and ll=318) then grbp<="010";
	end if;
	if (cc=89 and ll=318) then grbp<="010";
	end if;
	if (cc=114 and ll=318) then grbp<="010";
	end if;
	if (ll=318 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (ll=318 and cc>=122 and cc<137) then grbp<="010";
	end if;
	if (cc=148 and ll=318) then grbp<="010";
	end if;
	if (ll=318 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (cc=171 and ll=318) then grbp<="010";
	end if;
	if (ll=318 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=318) then grbp<="010";
	end if;
	if (cc=188 and ll=318) then grbp<="010";
	end if;
	if (ll=318 and cc>=188 and cc<197) then grbp<="010";
	end if;
	if (cc=210 and ll=318) then grbp<="010";
	end if;
	if (ll=318 and cc>=210 and cc<221) then grbp<="010";
	end if;
	if (ll=318 and cc>=246 and cc<249) then grbp<="010";
	end if;
	if (ll=319 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=319 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=37 and ll=319) then grbp<="010";
	end if;
	if (ll=319 and cc>=37 and cc<39) then grbp<="010";
	end if;
	if (cc=58 and ll=319) then grbp<="010";
	end if;
	if (cc=77 and ll=319) then grbp<="010";
	end if;
	if (cc=89 and ll=319) then grbp<="010";
	end if;
	if (cc=114 and ll=319) then grbp<="010";
	end if;
	if (ll=319 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (ll=319 and cc>=123 and cc<140) then grbp<="010";
	end if;
	if (ll=319 and cc>=144 and cc<153) then grbp<="010";
	end if;
	if (ll=319 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=319) then grbp<="010";
	end if;
	if (cc=188 and ll=319) then grbp<="010";
	end if;
	if (ll=319 and cc>=188 and cc<198) then grbp<="010";
	end if;
	if (cc=211 and ll=319) then grbp<="010";
	end if;
	if (ll=319 and cc>=211 and cc<220) then grbp<="010";
	end if;
	if (ll=319 and cc>=245 and cc<247) then grbp<="010";
	end if;
	if (ll=320 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=320 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=37 and ll=320) then grbp<="010";
	end if;
	if (cc=42 and ll=320) then grbp<="010";
	end if;
	if (cc=63 and ll=320) then grbp<="010";
	end if;
	if (cc=89 and ll=320) then grbp<="010";
	end if;
	if (cc=93 and ll=320) then grbp<="010";
	end if;
	if (cc=114 and ll=320) then grbp<="010";
	end if;
	if (ll=320 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (ll=320 and cc>=124 and cc<140) then grbp<="010";
	end if;
	if (ll=320 and cc>=144 and cc<153) then grbp<="010";
	end if;
	if (ll=320 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=320) then grbp<="010";
	end if;
	if (cc=187 and ll=320) then grbp<="010";
	end if;
	if (ll=320 and cc>=187 and cc<200) then grbp<="010";
	end if;
	if (ll=320 and cc>=210 and cc<220) then grbp<="010";
	end if;
	if (ll=320 and cc>=243 and cc<246) then grbp<="010";
	end if;
	if (ll=321 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=321 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=321 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (cc=89 and ll=321) then grbp<="010";
	end if;
	if (cc=93 and ll=321) then grbp<="010";
	end if;
	if (cc=115 and ll=321) then grbp<="010";
	end if;
	if (ll=321 and cc>=115 and cc<118) then grbp<="010";
	end if;
	if (ll=321 and cc>=120 and cc<136) then grbp<="010";
	end if;
	if (ll=321 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=321 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=321) then grbp<="010";
	end if;
	if (cc=187 and ll=321) then grbp<="010";
	end if;
	if (ll=321 and cc>=187 and cc<204) then grbp<="010";
	end if;
	if (ll=321 and cc>=207 and cc<209) then grbp<="010";
	end if;
	if (ll=321 and cc>=210 and cc<220) then grbp<="010";
	end if;
	if (ll=321 and cc>=242 and cc<244) then grbp<="010";
	end if;
	if (ll=322 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=322 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=75 and ll=322) then grbp<="010";
	end if;
	if (cc=87 and ll=322) then grbp<="010";
	end if;
	if (cc=89 and ll=322) then grbp<="010";
	end if;
	if (cc=115 and ll=322) then grbp<="010";
	end if;
	if (ll=322 and cc>=115 and cc<132) then grbp<="010";
	end if;
	if (ll=322 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (cc=171 and ll=322) then grbp<="010";
	end if;
	if (ll=322 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=184 and ll=322) then grbp<="010";
	end if;
	if (cc=187 and ll=322) then grbp<="010";
	end if;
	if (ll=322 and cc>=187 and cc<204) then grbp<="010";
	end if;
	if (ll=322 and cc>=208 and cc<220) then grbp<="010";
	end if;
	if (ll=322 and cc>=241 and cc<243) then grbp<="010";
	end if;
	if (ll=323 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=323 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=37 and ll=323) then grbp<="010";
	end if;
	if (cc=76 and ll=323) then grbp<="010";
	end if;
	if (cc=87 and ll=323) then grbp<="010";
	end if;
	if (ll=323 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=323 and cc>=115 and cc<137) then grbp<="010";
	end if;
	if (cc=153 and ll=323) then grbp<="010";
	end if;
	if (cc=171 and ll=323) then grbp<="010";
	end if;
	if (ll=323 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (ll=323 and cc>=181 and cc<183) then grbp<="010";
	end if;
	if (cc=187 and ll=323) then grbp<="010";
	end if;
	if (ll=323 and cc>=187 and cc<207) then grbp<="010";
	end if;
	if (ll=323 and cc>=208 and cc<220) then grbp<="010";
	end if;
	if (ll=323 and cc>=240 and cc<242) then grbp<="010";
	end if;
	if (ll=324 and cc>=10 and cc<17) then grbp<="010";
	end if;
	if (ll=324 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (ll=324 and cc>=34 and cc<36) then grbp<="010";
	end if;
	if (ll=324 and cc>=37 and cc<39) then grbp<="010";
	end if;
	if (cc=80 and ll=324) then grbp<="010";
	end if;
	if (cc=87 and ll=324) then grbp<="010";
	end if;
	if (ll=324 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (cc=116 and ll=324) then grbp<="010";
	end if;
	if (ll=324 and cc>=116 and cc<138) then grbp<="010";
	end if;
	if (ll=324 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (cc=171 and ll=324) then grbp<="010";
	end if;
	if (ll=324 and cc>=171 and cc<183) then grbp<="010";
	end if;
	if (ll=324 and cc>=187 and cc<220) then grbp<="010";
	end if;
	if (ll=324 and cc>=240 and cc<242) then grbp<="010";
	end if;
	if (cc=11 and ll=325) then grbp<="010";
	end if;
	if (ll=325 and cc>=11 and cc<17) then grbp<="010";
	end if;
	if (ll=325 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=38 and ll=325) then grbp<="010";
	end if;
	if (cc=43 and ll=325) then grbp<="010";
	end if;
	if (cc=88 and ll=325) then grbp<="010";
	end if;
	if (cc=93 and ll=325) then grbp<="010";
	end if;
	if (cc=116 and ll=325) then grbp<="010";
	end if;
	if (ll=325 and cc>=116 and cc<138) then grbp<="010";
	end if;
	if (ll=325 and cc>=139 and cc<146) then grbp<="010";
	end if;
	if (ll=325 and cc>=171 and cc<182) then grbp<="010";
	end if;
	if (ll=325 and cc>=187 and cc<220) then grbp<="010";
	end if;
	if (ll=325 and cc>=240 and cc<242) then grbp<="010";
	end if;
	if (ll=325 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=326) then grbp<="010";
	end if;
	if (ll=326 and cc>=11 and cc<18) then grbp<="010";
	end if;
	if (ll=326 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=37 and ll=326) then grbp<="010";
	end if;
	if (cc=43 and ll=326) then grbp<="010";
	end if;
	if (cc=50 and ll=326) then grbp<="010";
	end if;
	if (cc=74 and ll=326) then grbp<="010";
	end if;
	if (cc=88 and ll=326) then grbp<="010";
	end if;
	if (cc=93 and ll=326) then grbp<="010";
	end if;
	if (cc=116 and ll=326) then grbp<="010";
	end if;
	if (ll=326 and cc>=116 and cc<146) then grbp<="010";
	end if;
	if (ll=326 and cc>=170 and cc<182) then grbp<="010";
	end if;
	if (cc=187 and ll=326) then grbp<="010";
	end if;
	if (ll=326 and cc>=187 and cc<220) then grbp<="010";
	end if;
	if (ll=326 and cc>=239 and cc<241) then grbp<="010";
	end if;
	if (ll=326 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=327) then grbp<="010";
	end if;
	if (ll=327 and cc>=11 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=327) then grbp<="010";
	end if;
	if (cc=34 and ll=327) then grbp<="010";
	end if;
	if (cc=43 and ll=327) then grbp<="010";
	end if;
	if (cc=59 and ll=327) then grbp<="010";
	end if;
	if (cc=74 and ll=327) then grbp<="010";
	end if;
	if (ll=327 and cc>=74 and cc<76) then grbp<="010";
	end if;
	if (cc=93 and ll=327) then grbp<="010";
	end if;
	if (cc=116 and ll=327) then grbp<="010";
	end if;
	if (ll=327 and cc>=116 and cc<146) then grbp<="010";
	end if;
	if (ll=327 and cc>=171 and cc<183) then grbp<="010";
	end if;
	if (ll=327 and cc>=185 and cc<220) then grbp<="010";
	end if;
	if (ll=327 and cc>=239 and cc<241) then grbp<="010";
	end if;
	if (ll=327 and cc>=247 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=328) then grbp<="010";
	end if;
	if (cc=13 and ll=328) then grbp<="010";
	end if;
	if (ll=328 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (cc=34 and ll=328) then grbp<="010";
	end if;
	if (cc=43 and ll=328) then grbp<="010";
	end if;
	if (cc=51 and ll=328) then grbp<="010";
	end if;
	if (cc=80 and ll=328) then grbp<="010";
	end if;
	if (cc=88 and ll=328) then grbp<="010";
	end if;
	if (cc=93 and ll=328) then grbp<="010";
	end if;
	if (cc=116 and ll=328) then grbp<="010";
	end if;
	if (ll=328 and cc>=116 and cc<146) then grbp<="010";
	end if;
	if (cc=171 and ll=328) then grbp<="010";
	end if;
	if (ll=328 and cc>=171 and cc<183) then grbp<="010";
	end if;
	if (ll=328 and cc>=185 and cc<220) then grbp<="010";
	end if;
	if (ll=328 and cc>=238 and cc<240) then grbp<="010";
	end if;
	if (ll=328 and cc>=246 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=329) then grbp<="010";
	end if;
	if (ll=329 and cc>=0 and cc<3) then grbp<="010";
	end if;
	if (ll=329 and cc>=13 and cc<18) then grbp<="010";
	end if;
	if (ll=329 and cc>=31 and cc<33) then grbp<="010";
	end if;
	if (cc=51 and ll=329) then grbp<="010";
	end if;
	if (cc=80 and ll=329) then grbp<="010";
	end if;
	if (cc=88 and ll=329) then grbp<="010";
	end if;
	if (cc=93 and ll=329) then grbp<="010";
	end if;
	if (cc=116 and ll=329) then grbp<="010";
	end if;
	if (ll=329 and cc>=116 and cc<146) then grbp<="010";
	end if;
	if (cc=171 and ll=329) then grbp<="010";
	end if;
	if (ll=329 and cc>=171 and cc<181) then grbp<="010";
	end if;
	if (ll=329 and cc>=186 and cc<220) then grbp<="010";
	end if;
	if (ll=329 and cc>=237 and cc<239) then grbp<="010";
	end if;
	if (ll=329 and cc>=246 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=330) then grbp<="010";
	end if;
	if (ll=330 and cc>=0 and cc<4) then grbp<="010";
	end if;
	if (ll=330 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=330 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (ll=330 and cc>=34 and cc<36) then grbp<="010";
	end if;
	if (cc=51 and ll=330) then grbp<="010";
	end if;
	if (cc=60 and ll=330) then grbp<="010";
	end if;
	if (cc=80 and ll=330) then grbp<="010";
	end if;
	if (cc=88 and ll=330) then grbp<="010";
	end if;
	if (cc=93 and ll=330) then grbp<="010";
	end if;
	if (cc=116 and ll=330) then grbp<="010";
	end if;
	if (ll=330 and cc>=116 and cc<146) then grbp<="010";
	end if;
	if (ll=330 and cc>=171 and cc<182) then grbp<="010";
	end if;
	if (cc=186 and ll=330) then grbp<="010";
	end if;
	if (ll=330 and cc>=186 and cc<220) then grbp<="010";
	end if;
	if (cc=245 and ll=330) then grbp<="010";
	end if;
	if (ll=330 and cc>=245 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=331) then grbp<="010";
	end if;
	if (ll=331 and cc>=0 and cc<6) then grbp<="010";
	end if;
	if (ll=331 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=331 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=51 and ll=331) then grbp<="010";
	end if;
	if (cc=79 and ll=331) then grbp<="010";
	end if;
	if (ll=331 and cc>=79 and cc<81) then grbp<="010";
	end if;
	if (cc=88 and ll=331) then grbp<="010";
	end if;
	if (cc=93 and ll=331) then grbp<="010";
	end if;
	if (cc=116 and ll=331) then grbp<="010";
	end if;
	if (ll=331 and cc>=116 and cc<145) then grbp<="010";
	end if;
	if (ll=331 and cc>=171 and cc<180) then grbp<="010";
	end if;
	if (cc=183 and ll=331) then grbp<="010";
	end if;
	if (cc=186 and ll=331) then grbp<="010";
	end if;
	if (ll=331 and cc>=186 and cc<220) then grbp<="010";
	end if;
	if (ll=331 and cc>=236 and cc<238) then grbp<="010";
	end if;
	if (ll=331 and cc>=245 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=332) then grbp<="010";
	end if;
	if (ll=332 and cc>=0 and cc<6) then grbp<="010";
	end if;
	if (cc=14 and ll=332) then grbp<="010";
	end if;
	if (ll=332 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=332 and cc>=30 and cc<35) then grbp<="010";
	end if;
	if (cc=45 and ll=332) then grbp<="010";
	end if;
	if (ll=332 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=77 and ll=332) then grbp<="010";
	end if;
	if (cc=79 and ll=332) then grbp<="010";
	end if;
	if (cc=88 and ll=332) then grbp<="010";
	end if;
	if (cc=93 and ll=332) then grbp<="010";
	end if;
	if (cc=116 and ll=332) then grbp<="010";
	end if;
	if (ll=332 and cc>=116 and cc<145) then grbp<="010";
	end if;
	if (ll=332 and cc>=171 and cc<174) then grbp<="010";
	end if;
	if (ll=332 and cc>=175 and cc<184) then grbp<="010";
	end if;
	if (ll=332 and cc>=185 and cc<220) then grbp<="010";
	end if;
	if (cc=242 and ll=332) then grbp<="010";
	end if;
	if (ll=332 and cc>=242 and cc<251) then grbp<="010";
	end if;
	if (cc=2 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=2 and cc<7) then grbp<="010";
	end if;
	if (cc=14 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=333 and cc>=29 and cc<35) then grbp<="010";
	end if;
	if (ll=333 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=54 and ll=333) then grbp<="010";
	end if;
	if (cc=59 and ll=333) then grbp<="010";
	end if;
	if (cc=80 and ll=333) then grbp<="010";
	end if;
	if (cc=83 and ll=333) then grbp<="010";
	end if;
	if (cc=87 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=87 and cc<89) then grbp<="010";
	end if;
	if (cc=117 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=117 and cc<144) then grbp<="010";
	end if;
	if (cc=172 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (cc=177 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=177 and cc<182) then grbp<="010";
	end if;
	if (cc=185 and ll=333) then grbp<="010";
	end if;
	if (ll=333 and cc>=185 and cc<220) then grbp<="010";
	end if;
	if (ll=333 and cc>=235 and cc<237) then grbp<="010";
	end if;
	if (ll=333 and cc>=240 and cc<251) then grbp<="010";
	end if;
	if (cc=3 and ll=334) then grbp<="010";
	end if;
	if (ll=334 and cc>=3 and cc<10) then grbp<="010";
	end if;
	if (ll=334 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=334 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=45 and ll=334) then grbp<="010";
	end if;
	if (ll=334 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=78 and ll=334) then grbp<="010";
	end if;
	if (cc=80 and ll=334) then grbp<="010";
	end if;
	if (cc=83 and ll=334) then grbp<="010";
	end if;
	if (cc=88 and ll=334) then grbp<="010";
	end if;
	if (cc=117 and ll=334) then grbp<="010";
	end if;
	if (ll=334 and cc>=117 and cc<144) then grbp<="010";
	end if;
	if (cc=172 and ll=334) then grbp<="010";
	end if;
	if (ll=334 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=334 and cc>=177 and cc<180) then grbp<="010";
	end if;
	if (cc=185 and ll=334) then grbp<="010";
	end if;
	if (ll=334 and cc>=185 and cc<189) then grbp<="010";
	end if;
	if (ll=334 and cc>=190 and cc<220) then grbp<="010";
	end if;
	if (ll=334 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (ll=334 and cc>=240 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=335) then grbp<="010";
	end if;
	if (ll=335 and cc>=4 and cc<11) then grbp<="010";
	end if;
	if (ll=335 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=335 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (cc=45 and ll=335) then grbp<="010";
	end if;
	if (ll=335 and cc>=45 and cc<47) then grbp<="010";
	end if;
	if (cc=65 and ll=335) then grbp<="010";
	end if;
	if (cc=73 and ll=335) then grbp<="010";
	end if;
	if (cc=78 and ll=335) then grbp<="010";
	end if;
	if (ll=335 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (cc=87 and ll=335) then grbp<="010";
	end if;
	if (cc=112 and ll=335) then grbp<="010";
	end if;
	if (cc=117 and ll=335) then grbp<="010";
	end if;
	if (ll=335 and cc>=117 and cc<144) then grbp<="010";
	end if;
	if (ll=335 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=335 and cc>=177 and cc<180) then grbp<="010";
	end if;
	if (cc=185 and ll=335) then grbp<="010";
	end if;
	if (ll=335 and cc>=185 and cc<220) then grbp<="010";
	end if;
	if (ll=335 and cc>=233 and cc<235) then grbp<="010";
	end if;
	if (ll=335 and cc>=238 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=336) then grbp<="010";
	end if;
	if (ll=336 and cc>=5 and cc<11) then grbp<="010";
	end if;
	if (ll=336 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=336 and cc>=29 and cc<33) then grbp<="010";
	end if;
	if (ll=336 and cc>=34 and cc<36) then grbp<="010";
	end if;
	if (cc=78 and ll=336) then grbp<="010";
	end if;
	if (ll=336 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (ll=336 and cc>=84 and cc<86) then grbp<="010";
	end if;
	if (cc=111 and ll=336) then grbp<="010";
	end if;
	if (ll=336 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=336 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (ll=336 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=336 and cc>=177 and cc<180) then grbp<="010";
	end if;
	if (cc=185 and ll=336) then grbp<="010";
	end if;
	if (ll=336 and cc>=185 and cc<191) then grbp<="010";
	end if;
	if (ll=336 and cc>=192 and cc<220) then grbp<="010";
	end if;
	if (cc=238 and ll=336) then grbp<="010";
	end if;
	if (ll=336 and cc>=238 and cc<251) then grbp<="010";
	end if;
	if (cc=6 and ll=337) then grbp<="010";
	end if;
	if (ll=337 and cc>=6 and cc<11) then grbp<="010";
	end if;
	if (ll=337 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=337 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=337 and cc>=33 and cc<36) then grbp<="010";
	end if;
	if (cc=51 and ll=337) then grbp<="010";
	end if;
	if (cc=84 and ll=337) then grbp<="010";
	end if;
	if (cc=93 and ll=337) then grbp<="010";
	end if;
	if (cc=111 and ll=337) then grbp<="010";
	end if;
	if (ll=337 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=337 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (ll=337 and cc>=172 and cc<174) then grbp<="010";
	end if;
	if (ll=337 and cc>=178 and cc<181) then grbp<="010";
	end if;
	if (cc=185 and ll=337) then grbp<="010";
	end if;
	if (ll=337 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=337 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=337 and cc>=191 and cc<220) then grbp<="010";
	end if;
	if (ll=337 and cc>=232 and cc<234) then grbp<="010";
	end if;
	if (ll=337 and cc>=237 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=338) then grbp<="010";
	end if;
	if (ll=338 and cc>=7 and cc<11) then grbp<="010";
	end if;
	if (ll=338 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=338 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=338 and cc>=33 and cc<36) then grbp<="010";
	end if;
	if (cc=50 and ll=338) then grbp<="010";
	end if;
	if (cc=84 and ll=338) then grbp<="010";
	end if;
	if (cc=93 and ll=338) then grbp<="010";
	end if;
	if (cc=111 and ll=338) then grbp<="010";
	end if;
	if (ll=338 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=338 and cc>=117 and cc<142) then grbp<="010";
	end if;
	if (cc=178 and ll=338) then grbp<="010";
	end if;
	if (cc=180 and ll=338) then grbp<="010";
	end if;
	if (cc=183 and ll=338) then grbp<="010";
	end if;
	if (cc=185 and ll=338) then grbp<="010";
	end if;
	if (ll=338 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (ll=338 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=338 and cc>=191 and cc<219) then grbp<="010";
	end if;
	if (ll=338 and cc>=232 and cc<234) then grbp<="010";
	end if;
	if (ll=338 and cc>=237 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=339) then grbp<="010";
	end if;
	if (ll=339 and cc>=7 and cc<11) then grbp<="010";
	end if;
	if (ll=339 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=339 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=339 and cc>=33 and cc<36) then grbp<="010";
	end if;
	if (ll=339 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (cc=93 and ll=339) then grbp<="010";
	end if;
	if (cc=111 and ll=339) then grbp<="010";
	end if;
	if (ll=339 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=339 and cc>=117 and cc<142) then grbp<="010";
	end if;
	if (cc=183 and ll=339) then grbp<="010";
	end if;
	if (cc=185 and ll=339) then grbp<="010";
	end if;
	if (ll=339 and cc>=185 and cc<187) then grbp<="010";
	end if;
	if (cc=190 and ll=339) then grbp<="010";
	end if;
	if (ll=339 and cc>=190 and cc<219) then grbp<="010";
	end if;
	if (cc=236 and ll=339) then grbp<="010";
	end if;
	if (ll=339 and cc>=236 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=340) then grbp<="010";
	end if;
	if (cc=8 and ll=340) then grbp<="010";
	end if;
	if (ll=340 and cc>=8 and cc<11) then grbp<="010";
	end if;
	if (ll=340 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=340 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=340 and cc>=33 and cc<35) then grbp<="010";
	end if;
	if (cc=81 and ll=340) then grbp<="010";
	end if;
	if (cc=85 and ll=340) then grbp<="010";
	end if;
	if (cc=93 and ll=340) then grbp<="010";
	end if;
	if (cc=111 and ll=340) then grbp<="010";
	end if;
	if (ll=340 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=340 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (cc=173 and ll=340) then grbp<="010";
	end if;
	if (cc=178 and ll=340) then grbp<="010";
	end if;
	if (cc=183 and ll=340) then grbp<="010";
	end if;
	if (ll=340 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (cc=190 and ll=340) then grbp<="010";
	end if;
	if (ll=340 and cc>=190 and cc<194) then grbp<="010";
	end if;
	if (ll=340 and cc>=195 and cc<219) then grbp<="010";
	end if;
	if (cc=236 and ll=340) then grbp<="010";
	end if;
	if (ll=340 and cc>=236 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=341) then grbp<="010";
	end if;
	if (cc=9 and ll=341) then grbp<="010";
	end if;
	if (ll=341 and cc>=9 and cc<11) then grbp<="010";
	end if;
	if (ll=341 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=341 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=108 and ll=341) then grbp<="010";
	end if;
	if (cc=111 and ll=341) then grbp<="010";
	end if;
	if (ll=341 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=341 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (ll=341 and cc>=177 and cc<180) then grbp<="010";
	end if;
	if (ll=341 and cc>=183 and cc<187) then grbp<="010";
	end if;
	if (ll=341 and cc>=190 and cc<194) then grbp<="010";
	end if;
	if (ll=341 and cc>=195 and cc<219) then grbp<="010";
	end if;
	if (cc=235 and ll=341) then grbp<="010";
	end if;
	if (ll=341 and cc>=235 and cc<251) then grbp<="010";
	end if;
	if (cc=1 and ll=342) then grbp<="010";
	end if;
	if (cc=9 and ll=342) then grbp<="010";
	end if;
	if (ll=342 and cc>=9 and cc<12) then grbp<="010";
	end if;
	if (ll=342 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=342 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=108 and ll=342) then grbp<="010";
	end if;
	if (cc=111 and ll=342) then grbp<="010";
	end if;
	if (ll=342 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=342 and cc>=117 and cc<142) then grbp<="010";
	end if;
	if (cc=178 and ll=342) then grbp<="010";
	end if;
	if (cc=180 and ll=342) then grbp<="010";
	end if;
	if (cc=184 and ll=342) then grbp<="010";
	end if;
	if (ll=342 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (cc=192 and ll=342) then grbp<="010";
	end if;
	if (ll=342 and cc>=192 and cc<219) then grbp<="010";
	end if;
	if (ll=342 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=342 and cc>=235 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=343) then grbp<="010";
	end if;
	if (ll=343 and cc>=0 and cc<2) then grbp<="010";
	end if;
	if (ll=343 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=343 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=343 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=343 and cc>=32 and cc<34) then grbp<="010";
	end if;
	if (cc=84 and ll=343) then grbp<="010";
	end if;
	if (cc=108 and ll=343) then grbp<="010";
	end if;
	if (cc=111 and ll=343) then grbp<="010";
	end if;
	if (ll=343 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=343 and cc>=117 and cc<142) then grbp<="010";
	end if;
	if (cc=184 and ll=343) then grbp<="010";
	end if;
	if (ll=343 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=343 and cc>=193 and cc<219) then grbp<="010";
	end if;
	if (ll=343 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=343 and cc>=235 and cc<251) then grbp<="010";
	end if;
	if (cc=0 and ll=344) then grbp<="010";
	end if;
	if (ll=344 and cc>=0 and cc<3) then grbp<="010";
	end if;
	if (ll=344 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=344 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=344 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=63 and ll=344) then grbp<="010";
	end if;
	if (cc=81 and ll=344) then grbp<="010";
	end if;
	if (ll=344 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (cc=111 and ll=344) then grbp<="010";
	end if;
	if (ll=344 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=344 and cc>=117 and cc<142) then grbp<="010";
	end if;
	if (cc=177 and ll=344) then grbp<="010";
	end if;
	if (cc=184 and ll=344) then grbp<="010";
	end if;
	if (ll=344 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (cc=192 and ll=344) then grbp<="010";
	end if;
	if (ll=344 and cc>=192 and cc<218) then grbp<="010";
	end if;
	if (ll=344 and cc>=231 and cc<233) then grbp<="010";
	end if;
	if (ll=344 and cc>=234 and cc<251) then grbp<="010";
	end if;
	if (cc=1 and ll=345) then grbp<="010";
	end if;
	if (ll=345 and cc>=1 and cc<3) then grbp<="010";
	end if;
	if (ll=345 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=345 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=345 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=34 and ll=345) then grbp<="010";
	end if;
	if (cc=52 and ll=345) then grbp<="010";
	end if;
	if (cc=58 and ll=345) then grbp<="010";
	end if;
	if (cc=73 and ll=345) then grbp<="010";
	end if;
	if (cc=81 and ll=345) then grbp<="010";
	end if;
	if (ll=345 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (cc=111 and ll=345) then grbp<="010";
	end if;
	if (ll=345 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=345 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (ll=345 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=345 and cc>=192 and cc<218) then grbp<="010";
	end if;
	if (ll=345 and cc>=230 and cc<232) then grbp<="010";
	end if;
	if (ll=345 and cc>=234 and cc<251) then grbp<="010";
	end if;
	if (cc=2 and ll=346) then grbp<="010";
	end if;
	if (cc=10 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=346 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=346 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=346 and cc>=32 and cc<34) then grbp<="010";
	end if;
	if (cc=63 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (ll=346 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (cc=111 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=346 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (cc=184 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=346 and cc>=187 and cc<191) then grbp<="010";
	end if;
	if (ll=346 and cc>=192 and cc<199) then grbp<="010";
	end if;
	if (ll=346 and cc>=200 and cc<218) then grbp<="010";
	end if;
	if (ll=346 and cc>=230 and cc<232) then grbp<="010";
	end if;
	if (ll=346 and cc>=233 and cc<251) then grbp<="010";
	end if;
	if (cc=2 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=2 and cc<4) then grbp<="010";
	end if;
	if (ll=347 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=347 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=32 and cc<34) then grbp<="010";
	end if;
	if (ll=347 and cc>=51 and cc<53) then grbp<="010";
	end if;
	if (cc=86 and ll=347) then grbp<="010";
	end if;
	if (cc=111 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=347 and cc>=117 and cc<143) then grbp<="010";
	end if;
	if (cc=184 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=184 and cc<189) then grbp<="010";
	end if;
	if (ll=347 and cc>=191 and cc<195) then grbp<="010";
	end if;
	if (ll=347 and cc>=196 and cc<218) then grbp<="010";
	end if;
	if (ll=347 and cc>=230 and cc<251) then grbp<="010";
	end if;
	if (cc=2 and ll=348) then grbp<="010";
	end if;
	if (ll=348 and cc>=2 and cc<4) then grbp<="010";
	end if;
	if (ll=348 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=348 and cc>=14 and cc<18) then grbp<="010";
	end if;
	if (ll=348 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=348 and cc>=32 and cc<35) then grbp<="010";
	end if;
	if (cc=75 and ll=348) then grbp<="010";
	end if;
	if (cc=84 and ll=348) then grbp<="010";
	end if;
	if (cc=110 and ll=348) then grbp<="010";
	end if;
	if (ll=348 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=348 and cc>=117 and cc<144) then grbp<="010";
	end if;
	if (cc=184 and ll=348) then grbp<="010";
	end if;
	if (ll=348 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=348 and cc>=188 and cc<218) then grbp<="010";
	end if;
	if (ll=348 and cc>=229 and cc<251) then grbp<="010";
	end if;
	if (cc=3 and ll=349) then grbp<="010";
	end if;
	if (cc=10 and ll=349) then grbp<="010";
	end if;
	if (ll=349 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=349 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=349 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (ll=349 and cc>=32 and cc<35) then grbp<="010";
	end if;
	if (cc=52 and ll=349) then grbp<="010";
	end if;
	if (cc=59 and ll=349) then grbp<="010";
	end if;
	if (cc=65 and ll=349) then grbp<="010";
	end if;
	if (cc=75 and ll=349) then grbp<="010";
	end if;
	if (cc=86 and ll=349) then grbp<="010";
	end if;
	if (cc=110 and ll=349) then grbp<="010";
	end if;
	if (ll=349 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=349 and cc>=118 and cc<143) then grbp<="010";
	end if;
	if (cc=182 and ll=349) then grbp<="010";
	end if;
	if (cc=184 and ll=349) then grbp<="010";
	end if;
	if (ll=349 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=349 and cc>=189 and cc<217) then grbp<="010";
	end if;
	if (ll=349 and cc>=229 and cc<251) then grbp<="010";
	end if;
	if (cc=3 and ll=350) then grbp<="010";
	end if;
	if (cc=10 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=10 and cc<12) then grbp<="010";
	end if;
	if (ll=350 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=350 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (ll=350 and cc>=33 and cc<35) then grbp<="010";
	end if;
	if (cc=60 and ll=350) then grbp<="010";
	end if;
	if (cc=75 and ll=350) then grbp<="010";
	end if;
	if (cc=110 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=350 and cc>=118 and cc<144) then grbp<="010";
	end if;
	if (cc=184 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=350 and cc>=188 and cc<215) then grbp<="010";
	end if;
	if (ll=350 and cc>=229 and cc<251) then grbp<="010";
	end if;
	if (cc=3 and ll=351) then grbp<="010";
	end if;
	if (cc=11 and ll=351) then grbp<="010";
	end if;
	if (cc=15 and ll=351) then grbp<="010";
	end if;
	if (ll=351 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=351 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (ll=351 and cc>=33 and cc<35) then grbp<="010";
	end if;
	if (cc=60 and ll=351) then grbp<="010";
	end if;
	if (cc=81 and ll=351) then grbp<="010";
	end if;
	if (cc=86 and ll=351) then grbp<="010";
	end if;
	if (cc=95 and ll=351) then grbp<="010";
	end if;
	if (cc=110 and ll=351) then grbp<="010";
	end if;
	if (ll=351 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=351 and cc>=118 and cc<144) then grbp<="010";
	end if;
	if (cc=184 and ll=351) then grbp<="010";
	end if;
	if (ll=351 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=351 and cc>=187 and cc<189) then grbp<="010";
	end if;
	if (ll=351 and cc>=190 and cc<214) then grbp<="010";
	end if;
	if (ll=351 and cc>=229 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=352) then grbp<="010";
	end if;
	if (cc=15 and ll=352) then grbp<="010";
	end if;
	if (ll=352 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=352 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=61 and ll=352) then grbp<="010";
	end if;
	if (cc=95 and ll=352) then grbp<="010";
	end if;
	if (cc=110 and ll=352) then grbp<="010";
	end if;
	if (ll=352 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=352 and cc>=118 and cc<145) then grbp<="010";
	end if;
	if (cc=184 and ll=352) then grbp<="010";
	end if;
	if (ll=352 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=352 and cc>=188 and cc<194) then grbp<="010";
	end if;
	if (ll=352 and cc>=195 and cc<214) then grbp<="010";
	end if;
	if (ll=352 and cc>=229 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=353) then grbp<="010";
	end if;
	if (cc=15 and ll=353) then grbp<="010";
	end if;
	if (ll=353 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=353 and cc>=29 and cc<34) then grbp<="010";
	end if;
	if (cc=85 and ll=353) then grbp<="010";
	end if;
	if (cc=95 and ll=353) then grbp<="010";
	end if;
	if (cc=110 and ll=353) then grbp<="010";
	end if;
	if (ll=353 and cc>=110 and cc<115) then grbp<="010";
	end if;
	if (ll=353 and cc>=118 and cc<145) then grbp<="010";
	end if;
	if (cc=182 and ll=353) then grbp<="010";
	end if;
	if (cc=184 and ll=353) then grbp<="010";
	end if;
	if (ll=353 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (ll=353 and cc>=188 and cc<191) then grbp<="010";
	end if;
	if (ll=353 and cc>=192 and cc<213) then grbp<="010";
	end if;
	if (ll=353 and cc>=228 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=354) then grbp<="010";
	end if;
	if (cc=11 and ll=354) then grbp<="010";
	end if;
	if (cc=15 and ll=354) then grbp<="010";
	end if;
	if (ll=354 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=354 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=85 and ll=354) then grbp<="010";
	end if;
	if (cc=95 and ll=354) then grbp<="010";
	end if;
	if (cc=109 and ll=354) then grbp<="010";
	end if;
	if (ll=354 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=354 and cc>=118 and cc<144) then grbp<="010";
	end if;
	if (ll=354 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=354 and cc>=188 and cc<213) then grbp<="010";
	end if;
	if (ll=354 and cc>=228 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=355) then grbp<="010";
	end if;
	if (cc=11 and ll=355) then grbp<="010";
	end if;
	if (cc=15 and ll=355) then grbp<="010";
	end if;
	if (ll=355 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=355 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=85 and ll=355) then grbp<="010";
	end if;
	if (cc=92 and ll=355) then grbp<="010";
	end if;
	if (cc=95 and ll=355) then grbp<="010";
	end if;
	if (cc=109 and ll=355) then grbp<="010";
	end if;
	if (ll=355 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=355 and cc>=118 and cc<144) then grbp<="010";
	end if;
	if (cc=184 and ll=355) then grbp<="010";
	end if;
	if (ll=355 and cc>=184 and cc<186) then grbp<="010";
	end if;
	if (cc=192 and ll=355) then grbp<="010";
	end if;
	if (ll=355 and cc>=192 and cc<212) then grbp<="010";
	end if;
	if (ll=355 and cc>=228 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=356) then grbp<="010";
	end if;
	if (cc=11 and ll=356) then grbp<="010";
	end if;
	if (cc=15 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=356 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=55 and ll=356) then grbp<="010";
	end if;
	if (cc=69 and ll=356) then grbp<="010";
	end if;
	if (cc=85 and ll=356) then grbp<="010";
	end if;
	if (cc=92 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=92 and cc<94) then grbp<="010";
	end if;
	if (cc=109 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=356 and cc>=118 and cc<144) then grbp<="010";
	end if;
	if (cc=176 and ll=356) then grbp<="010";
	end if;
	if (cc=182 and ll=356) then grbp<="010";
	end if;
	if (cc=184 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=184 and cc<187) then grbp<="010";
	end if;
	if (ll=356 and cc>=190 and cc<192) then grbp<="010";
	end if;
	if (ll=356 and cc>=193 and cc<212) then grbp<="010";
	end if;
	if (ll=356 and cc>=228 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=357) then grbp<="010";
	end if;
	if (cc=11 and ll=357) then grbp<="010";
	end if;
	if (cc=15 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=357 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=92 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=92 and cc<94) then grbp<="010";
	end if;
	if (cc=109 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=357 and cc>=118 and cc<146) then grbp<="010";
	end if;
	if (cc=182 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (cc=192 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=192 and cc<211) then grbp<="010";
	end if;
	if (ll=357 and cc>=227 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=358) then grbp<="010";
	end if;
	if (cc=11 and ll=358) then grbp<="010";
	end if;
	if (cc=15 and ll=358) then grbp<="010";
	end if;
	if (ll=358 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=358 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=85 and ll=358) then grbp<="010";
	end if;
	if (cc=87 and ll=358) then grbp<="010";
	end if;
	if (cc=92 and ll=358) then grbp<="010";
	end if;
	if (cc=95 and ll=358) then grbp<="010";
	end if;
	if (cc=109 and ll=358) then grbp<="010";
	end if;
	if (ll=358 and cc>=109 and cc<116) then grbp<="010";
	end if;
	if (ll=358 and cc>=117 and cc<146) then grbp<="010";
	end if;
	if (ll=358 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (cc=190 and ll=358) then grbp<="010";
	end if;
	if (ll=358 and cc>=190 and cc<192) then grbp<="010";
	end if;
	if (ll=358 and cc>=193 and cc<211) then grbp<="010";
	end if;
	if (ll=358 and cc>=227 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=359) then grbp<="010";
	end if;
	if (cc=11 and ll=359) then grbp<="010";
	end if;
	if (cc=15 and ll=359) then grbp<="010";
	end if;
	if (ll=359 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=359 and cc>=29 and cc<34) then grbp<="010";
	end if;
	if (cc=108 and ll=359) then grbp<="010";
	end if;
	if (ll=359 and cc>=108 and cc<116) then grbp<="010";
	end if;
	if (ll=359 and cc>=117 and cc<146) then grbp<="010";
	end if;
	if (ll=359 and cc>=182 and cc<185) then grbp<="010";
	end if;
	if (cc=190 and ll=359) then grbp<="010";
	end if;
	if (ll=359 and cc>=190 and cc<211) then grbp<="010";
	end if;
	if (ll=359 and cc>=227 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=360) then grbp<="010";
	end if;
	if (cc=11 and ll=360) then grbp<="010";
	end if;
	if (cc=15 and ll=360) then grbp<="010";
	end if;
	if (ll=360 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=360 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=108 and ll=360) then grbp<="010";
	end if;
	if (ll=360 and cc>=108 and cc<116) then grbp<="010";
	end if;
	if (ll=360 and cc>=117 and cc<146) then grbp<="010";
	end if;
	if (ll=360 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=360 and cc>=188 and cc<192) then grbp<="010";
	end if;
	if (ll=360 and cc>=193 and cc<211) then grbp<="010";
	end if;
	if (ll=360 and cc>=226 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=361) then grbp<="010";
	end if;
	if (cc=11 and ll=361) then grbp<="010";
	end if;
	if (cc=15 and ll=361) then grbp<="010";
	end if;
	if (ll=361 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=361 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (ll=361 and cc>=50 and cc<52) then grbp<="010";
	end if;
	if (cc=108 and ll=361) then grbp<="010";
	end if;
	if (ll=361 and cc>=108 and cc<116) then grbp<="010";
	end if;
	if (ll=361 and cc>=117 and cc<147) then grbp<="010";
	end if;
	if (cc=181 and ll=361) then grbp<="010";
	end if;
	if (ll=361 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=188 and ll=361) then grbp<="010";
	end if;
	if (ll=361 and cc>=188 and cc<192) then grbp<="010";
	end if;
	if (ll=361 and cc>=193 and cc<211) then grbp<="010";
	end if;
	if (ll=361 and cc>=226 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=362) then grbp<="010";
	end if;
	if (cc=11 and ll=362) then grbp<="010";
	end if;
	if (cc=15 and ll=362) then grbp<="010";
	end if;
	if (ll=362 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=362 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (ll=362 and cc>=50 and cc<52) then grbp<="010";
	end if;
	if (cc=92 and ll=362) then grbp<="010";
	end if;
	if (cc=107 and ll=362) then grbp<="010";
	end if;
	if (ll=362 and cc>=107 and cc<116) then grbp<="010";
	end if;
	if (ll=362 and cc>=117 and cc<145) then grbp<="010";
	end if;
	if (cc=181 and ll=362) then grbp<="010";
	end if;
	if (ll=362 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=188 and ll=362) then grbp<="010";
	end if;
	if (ll=362 and cc>=188 and cc<210) then grbp<="010";
	end if;
	if (ll=362 and cc>=226 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=363) then grbp<="010";
	end if;
	if (cc=11 and ll=363) then grbp<="010";
	end if;
	if (cc=15 and ll=363) then grbp<="010";
	end if;
	if (ll=363 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=363 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=107 and ll=363) then grbp<="010";
	end if;
	if (ll=363 and cc>=107 and cc<116) then grbp<="010";
	end if;
	if (ll=363 and cc>=117 and cc<145) then grbp<="010";
	end if;
	if (ll=363 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=189 and ll=363) then grbp<="010";
	end if;
	if (ll=363 and cc>=189 and cc<210) then grbp<="010";
	end if;
	if (ll=363 and cc>=226 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=364) then grbp<="010";
	end if;
	if (cc=11 and ll=364) then grbp<="010";
	end if;
	if (cc=15 and ll=364) then grbp<="010";
	end if;
	if (ll=364 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=364 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=79 and ll=364) then grbp<="010";
	end if;
	if (cc=106 and ll=364) then grbp<="010";
	end if;
	if (ll=364 and cc>=106 and cc<115) then grbp<="010";
	end if;
	if (ll=364 and cc>=117 and cc<147) then grbp<="010";
	end if;
	if (ll=364 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=364 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (ll=364 and cc>=191 and cc<210) then grbp<="010";
	end if;
	if (ll=364 and cc>=225 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=365) then grbp<="010";
	end if;
	if (cc=11 and ll=365) then grbp<="010";
	end if;
	if (cc=15 and ll=365) then grbp<="010";
	end if;
	if (ll=365 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=365 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=106 and ll=365) then grbp<="010";
	end if;
	if (ll=365 and cc>=106 and cc<115) then grbp<="010";
	end if;
	if (ll=365 and cc>=117 and cc<147) then grbp<="010";
	end if;
	if (ll=365 and cc>=181 and cc<186) then grbp<="010";
	end if;
	if (cc=190 and ll=365) then grbp<="010";
	end if;
	if (ll=365 and cc>=190 and cc<210) then grbp<="010";
	end if;
	if (ll=365 and cc>=225 and cc<251) then grbp<="010";
	end if;
	if (cc=4 and ll=366) then grbp<="010";
	end if;
	if (cc=11 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=366 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=366 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=105 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=105 and cc<115) then grbp<="010";
	end if;
	if (ll=366 and cc>=117 and cc<146) then grbp<="010";
	end if;
	if (ll=366 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=366 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (ll=366 and cc>=191 and cc<210) then grbp<="010";
	end if;
	if (ll=366 and cc>=225 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=367) then grbp<="010";
	end if;
	if (ll=367 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=367 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=367 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=50 and ll=367) then grbp<="010";
	end if;
	if (cc=80 and ll=367) then grbp<="010";
	end if;
	if (cc=89 and ll=367) then grbp<="010";
	end if;
	if (cc=91 and ll=367) then grbp<="010";
	end if;
	if (cc=97 and ll=367) then grbp<="010";
	end if;
	if (cc=105 and ll=367) then grbp<="010";
	end if;
	if (ll=367 and cc>=105 and cc<115) then grbp<="010";
	end if;
	if (ll=367 and cc>=117 and cc<148) then grbp<="010";
	end if;
	if (cc=181 and ll=367) then grbp<="010";
	end if;
	if (ll=367 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=367 and cc>=187 and cc<210) then grbp<="010";
	end if;
	if (ll=367 and cc>=224 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=368 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=368 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=79 and ll=368) then grbp<="010";
	end if;
	if (cc=84 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=84 and cc<88) then grbp<="010";
	end if;
	if (cc=96 and ll=368) then grbp<="010";
	end if;
	if (cc=105 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=105 and cc<115) then grbp<="010";
	end if;
	if (ll=368 and cc>=116 and cc<147) then grbp<="010";
	end if;
	if (cc=181 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=368 and cc>=187 and cc<210) then grbp<="010";
	end if;
	if (ll=368 and cc>=224 and cc<251) then grbp<="010";
	end if;
	if (cc=11 and ll=369) then grbp<="010";
	end if;
	if (ll=369 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=369 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=369 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=67 and ll=369) then grbp<="010";
	end if;
	if (cc=80 and ll=369) then grbp<="010";
	end if;
	if (cc=84 and ll=369) then grbp<="010";
	end if;
	if (cc=88 and ll=369) then grbp<="010";
	end if;
	if (cc=96 and ll=369) then grbp<="010";
	end if;
	if (cc=105 and ll=369) then grbp<="010";
	end if;
	if (ll=369 and cc>=105 and cc<115) then grbp<="010";
	end if;
	if (ll=369 and cc>=116 and cc<149) then grbp<="010";
	end if;
	if (ll=369 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=189 and ll=369) then grbp<="010";
	end if;
	if (ll=369 and cc>=189 and cc<210) then grbp<="010";
	end if;
	if (ll=369 and cc>=224 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=370) then grbp<="010";
	end if;
	if (cc=11 and ll=370) then grbp<="010";
	end if;
	if (ll=370 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=370 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=370 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=67 and ll=370) then grbp<="010";
	end if;
	if (cc=80 and ll=370) then grbp<="010";
	end if;
	if (cc=91 and ll=370) then grbp<="010";
	end if;
	if (cc=93 and ll=370) then grbp<="010";
	end if;
	if (cc=95 and ll=370) then grbp<="010";
	end if;
	if (ll=370 and cc>=95 and cc<97) then grbp<="010";
	end if;
	if (ll=370 and cc>=105 and cc<115) then grbp<="010";
	end if;
	if (ll=370 and cc>=116 and cc<149) then grbp<="010";
	end if;
	if (ll=370 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=370 and cc>=189 and cc<210) then grbp<="010";
	end if;
	if (ll=370 and cc>=224 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=371) then grbp<="010";
	end if;
	if (cc=12 and ll=371) then grbp<="010";
	end if;
	if (cc=15 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=371) then grbp<="010";
	end if;
	if (cc=80 and ll=371) then grbp<="010";
	end if;
	if (cc=87 and ll=371) then grbp<="010";
	end if;
	if (cc=93 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (cc=104 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=104 and cc<115) then grbp<="010";
	end if;
	if (ll=371 and cc>=116 and cc<148) then grbp<="010";
	end if;
	if (ll=371 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=190 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=190 and cc<210) then grbp<="010";
	end if;
	if (ll=371 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=372) then grbp<="010";
	end if;
	if (cc=12 and ll=372) then grbp<="010";
	end if;
	if (cc=15 and ll=372) then grbp<="010";
	end if;
	if (ll=372 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=372) then grbp<="010";
	end if;
	if (cc=67 and ll=372) then grbp<="010";
	end if;
	if (cc=84 and ll=372) then grbp<="010";
	end if;
	if (cc=96 and ll=372) then grbp<="010";
	end if;
	if (ll=372 and cc>=96 and cc<98) then grbp<="010";
	end if;
	if (ll=372 and cc>=104 and cc<115) then grbp<="010";
	end if;
	if (ll=372 and cc>=116 and cc<148) then grbp<="010";
	end if;
	if (ll=372 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=372 and cc>=188 and cc<210) then grbp<="010";
	end if;
	if (ll=372 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=373) then grbp<="010";
	end if;
	if (cc=11 and ll=373) then grbp<="010";
	end if;
	if (ll=373 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=373 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=373) then grbp<="010";
	end if;
	if (cc=82 and ll=373) then grbp<="010";
	end if;
	if (cc=84 and ll=373) then grbp<="010";
	end if;
	if (cc=97 and ll=373) then grbp<="010";
	end if;
	if (cc=104 and ll=373) then grbp<="010";
	end if;
	if (ll=373 and cc>=104 and cc<115) then grbp<="010";
	end if;
	if (ll=373 and cc>=116 and cc<148) then grbp<="010";
	end if;
	if (cc=181 and ll=373) then grbp<="010";
	end if;
	if (ll=373 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=373 and cc>=187 and cc<192) then grbp<="010";
	end if;
	if (ll=373 and cc>=193 and cc<210) then grbp<="010";
	end if;
	if (ll=373 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=374) then grbp<="010";
	end if;
	if (cc=11 and ll=374) then grbp<="010";
	end if;
	if (ll=374 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=374 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=374) then grbp<="010";
	end if;
	if (cc=75 and ll=374) then grbp<="010";
	end if;
	if (cc=104 and ll=374) then grbp<="010";
	end if;
	if (ll=374 and cc>=104 and cc<115) then grbp<="010";
	end if;
	if (ll=374 and cc>=116 and cc<150) then grbp<="010";
	end if;
	if (cc=181 and ll=374) then grbp<="010";
	end if;
	if (ll=374 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (cc=189 and ll=374) then grbp<="010";
	end if;
	if (ll=374 and cc>=189 and cc<210) then grbp<="010";
	end if;
	if (ll=374 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=375) then grbp<="010";
	end if;
	if (cc=12 and ll=375) then grbp<="010";
	end if;
	if (cc=15 and ll=375) then grbp<="010";
	end if;
	if (ll=375 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=375 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=104 and ll=375) then grbp<="010";
	end if;
	if (ll=375 and cc>=104 and cc<114) then grbp<="010";
	end if;
	if (ll=375 and cc>=116 and cc<148) then grbp<="010";
	end if;
	if (ll=375 and cc>=181 and cc<185) then grbp<="010";
	end if;
	if (ll=375 and cc>=187 and cc<211) then grbp<="010";
	end if;
	if (ll=375 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=376) then grbp<="010";
	end if;
	if (cc=12 and ll=376) then grbp<="010";
	end if;
	if (cc=15 and ll=376) then grbp<="010";
	end if;
	if (ll=376 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=376 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=44 and ll=376) then grbp<="010";
	end if;
	if (cc=66 and ll=376) then grbp<="010";
	end if;
	if (cc=69 and ll=376) then grbp<="010";
	end if;
	if (cc=78 and ll=376) then grbp<="010";
	end if;
	if (cc=103 and ll=376) then grbp<="010";
	end if;
	if (ll=376 and cc>=103 and cc<114) then grbp<="010";
	end if;
	if (ll=376 and cc>=115 and cc<150) then grbp<="010";
	end if;
	if (ll=376 and cc>=180 and cc<185) then grbp<="010";
	end if;
	if (cc=188 and ll=376) then grbp<="010";
	end if;
	if (ll=376 and cc>=188 and cc<190) then grbp<="010";
	end if;
	if (ll=376 and cc>=191 and cc<193) then grbp<="010";
	end if;
	if (ll=376 and cc>=194 and cc<211) then grbp<="010";
	end if;
	if (ll=376 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=377) then grbp<="010";
	end if;
	if (cc=11 and ll=377) then grbp<="010";
	end if;
	if (ll=377 and cc>=11 and cc<13) then grbp<="010";
	end if;
	if (ll=377 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=377) then grbp<="010";
	end if;
	if (cc=34 and ll=377) then grbp<="010";
	end if;
	if (cc=43 and ll=377) then grbp<="010";
	end if;
	if (cc=69 and ll=377) then grbp<="010";
	end if;
	if (cc=103 and ll=377) then grbp<="010";
	end if;
	if (ll=377 and cc>=103 and cc<114) then grbp<="010";
	end if;
	if (ll=377 and cc>=115 and cc<150) then grbp<="010";
	end if;
	if (ll=377 and cc>=180 and cc<191) then grbp<="010";
	end if;
	if (ll=377 and cc>=193 and cc<212) then grbp<="010";
	end if;
	if (ll=377 and cc>=223 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=378) then grbp<="010";
	end if;
	if (cc=12 and ll=378) then grbp<="010";
	end if;
	if (cc=15 and ll=378) then grbp<="010";
	end if;
	if (ll=378 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=378) then grbp<="010";
	end if;
	if (cc=34 and ll=378) then grbp<="010";
	end if;
	if (cc=85 and ll=378) then grbp<="010";
	end if;
	if (cc=103 and ll=378) then grbp<="010";
	end if;
	if (ll=378 and cc>=103 and cc<114) then grbp<="010";
	end if;
	if (ll=378 and cc>=115 and cc<150) then grbp<="010";
	end if;
	if (ll=378 and cc>=180 and cc<192) then grbp<="010";
	end if;
	if (ll=378 and cc>=195 and cc<213) then grbp<="010";
	end if;
	if (ll=378 and cc>=222 and cc<251) then grbp<="010";
	end if;
	if (cc=5 and ll=379) then grbp<="010";
	end if;
	if (cc=12 and ll=379) then grbp<="010";
	end if;
	if (cc=15 and ll=379) then grbp<="010";
	end if;
	if (ll=379 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (cc=32 and ll=379) then grbp<="010";
	end if;
	if (cc=34 and ll=379) then grbp<="010";
	end if;
	if (cc=65 and ll=379) then grbp<="010";
	end if;
	if (cc=70 and ll=379) then grbp<="010";
	end if;
	if (cc=103 and ll=379) then grbp<="010";
	end if;
	if (ll=379 and cc>=103 and cc<114) then grbp<="010";
	end if;
	if (ll=379 and cc>=115 and cc<151) then grbp<="010";
	end if;
	if (ll=379 and cc>=180 and cc<194) then grbp<="010";
	end if;
	if (cc=198 and ll=379) then grbp<="010";
	end if;
	if (ll=379 and cc>=198 and cc<214) then grbp<="010";
	end if;
	if (ll=379 and cc>=222 and cc<250) then grbp<="010";
	end if;
	if (cc=15 and ll=380) then grbp<="010";
	end if;
	if (ll=380 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=380 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=86 and ll=380) then grbp<="010";
	end if;
	if (cc=102 and ll=380) then grbp<="010";
	end if;
	if (ll=380 and cc>=102 and cc<113) then grbp<="010";
	end if;
	if (ll=380 and cc>=115 and cc<151) then grbp<="010";
	end if;
	if (ll=380 and cc>=181 and cc<196) then grbp<="010";
	end if;
	if (ll=380 and cc>=197 and cc<206) then grbp<="010";
	end if;
	if (ll=380 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=380 and cc>=222 and cc<250) then grbp<="010";
	end if;
	if (cc=12 and ll=381) then grbp<="010";
	end if;
	if (cc=15 and ll=381) then grbp<="010";
	end if;
	if (ll=381 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=381 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=102 and ll=381) then grbp<="010";
	end if;
	if (ll=381 and cc>=102 and cc<113) then grbp<="010";
	end if;
	if (ll=381 and cc>=115 and cc<152) then grbp<="010";
	end if;
	if (ll=381 and cc>=181 and cc<197) then grbp<="010";
	end if;
	if (ll=381 and cc>=198 and cc<207) then grbp<="010";
	end if;
	if (ll=381 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=381 and cc>=222 and cc<250) then grbp<="010";
	end if;
	if (cc=12 and ll=382) then grbp<="010";
	end if;
	if (cc=15 and ll=382) then grbp<="010";
	end if;
	if (ll=382 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=382 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=84 and ll=382) then grbp<="010";
	end if;
	if (cc=102 and ll=382) then grbp<="010";
	end if;
	if (ll=382 and cc>=102 and cc<113) then grbp<="010";
	end if;
	if (ll=382 and cc>=114 and cc<152) then grbp<="010";
	end if;
	if (ll=382 and cc>=181 and cc<206) then grbp<="010";
	end if;
	if (ll=382 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=382 and cc>=222 and cc<249) then grbp<="010";
	end if;
	if (cc=12 and ll=383) then grbp<="010";
	end if;
	if (cc=15 and ll=383) then grbp<="010";
	end if;
	if (ll=383 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=383 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (cc=78 and ll=383) then grbp<="010";
	end if;
	if (cc=102 and ll=383) then grbp<="010";
	end if;
	if (ll=383 and cc>=102 and cc<113) then grbp<="010";
	end if;
	if (ll=383 and cc>=114 and cc<150) then grbp<="010";
	end if;
	if (cc=181 and ll=383) then grbp<="010";
	end if;
	if (ll=383 and cc>=181 and cc<206) then grbp<="010";
	end if;
	if (ll=383 and cc>=208 and cc<214) then grbp<="010";
	end if;
	if (ll=383 and cc>=221 and cc<249) then grbp<="010";
	end if;
	if (cc=12 and ll=384) then grbp<="010";
	end if;
	if (cc=15 and ll=384) then grbp<="010";
	end if;
	if (ll=384 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=384 and cc>=30 and cc<35) then grbp<="010";
	end if;
	if (ll=384 and cc>=83 and cc<85) then grbp<="010";
	end if;
	if (ll=384 and cc>=101 and cc<112) then grbp<="010";
	end if;
	if (ll=384 and cc>=114 and cc<153) then grbp<="010";
	end if;
	if (ll=384 and cc>=181 and cc<184) then grbp<="010";
	end if;
	if (ll=384 and cc>=185 and cc<204) then grbp<="010";
	end if;
	if (ll=384 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=384 and cc>=221 and cc<249) then grbp<="010";
	end if;
	if (cc=12 and ll=385) then grbp<="010";
	end if;
	if (cc=15 and ll=385) then grbp<="010";
	end if;
	if (ll=385 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=385 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (cc=84 and ll=385) then grbp<="010";
	end if;
	if (ll=385 and cc>=84 and cc<86) then grbp<="010";
	end if;
	if (ll=385 and cc>=101 and cc<112) then grbp<="010";
	end if;
	if (ll=385 and cc>=114 and cc<151) then grbp<="010";
	end if;
	if (ll=385 and cc>=181 and cc<186) then grbp<="010";
	end if;
	if (ll=385 and cc>=187 and cc<205) then grbp<="010";
	end if;
	if (ll=385 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=385 and cc>=221 and cc<248) then grbp<="010";
	end if;
	if (ll=386 and cc>=12 and cc<14) then grbp<="010";
	end if;
	if (ll=386 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=386 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (cc=84 and ll=386) then grbp<="010";
	end if;
	if (cc=100 and ll=386) then grbp<="010";
	end if;
	if (ll=386 and cc>=100 and cc<112) then grbp<="010";
	end if;
	if (ll=386 and cc>=113 and cc<151) then grbp<="010";
	end if;
	if (ll=386 and cc>=182 and cc<205) then grbp<="010";
	end if;
	if (ll=386 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=386 and cc>=221 and cc<248) then grbp<="010";
	end if;
	if (ll=387 and cc>=12 and cc<14) then grbp<="010";
	end if;
	if (ll=387 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=387 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=100 and ll=387) then grbp<="010";
	end if;
	if (ll=387 and cc>=100 and cc<111) then grbp<="010";
	end if;
	if (ll=387 and cc>=113 and cc<152) then grbp<="010";
	end if;
	if (ll=387 and cc>=182 and cc<206) then grbp<="010";
	end if;
	if (cc=211 and ll=387) then grbp<="010";
	end if;
	if (ll=387 and cc>=211 and cc<213) then grbp<="010";
	end if;
	if (ll=387 and cc>=220 and cc<247) then grbp<="010";
	end if;
	if (ll=388 and cc>=12 and cc<14) then grbp<="010";
	end if;
	if (ll=388 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=388 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (cc=81 and ll=388) then grbp<="010";
	end if;
	if (cc=100 and ll=388) then grbp<="010";
	end if;
	if (ll=388 and cc>=100 and cc<111) then grbp<="010";
	end if;
	if (ll=388 and cc>=113 and cc<153) then grbp<="010";
	end if;
	if (ll=388 and cc>=182 and cc<194) then grbp<="010";
	end if;
	if (ll=388 and cc>=196 and cc<206) then grbp<="010";
	end if;
	if (cc=220 and ll=388) then grbp<="010";
	end if;
	if (ll=388 and cc>=220 and cc<247) then grbp<="010";
	end if;
	if (cc=15 and ll=389) then grbp<="010";
	end if;
	if (ll=389 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=389 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (cc=100 and ll=389) then grbp<="010";
	end if;
	if (ll=389 and cc>=100 and cc<110) then grbp<="010";
	end if;
	if (ll=389 and cc>=113 and cc<153) then grbp<="010";
	end if;
	if (ll=389 and cc>=182 and cc<194) then grbp<="010";
	end if;
	if (ll=389 and cc>=202 and cc<208) then grbp<="010";
	end if;
	if (ll=389 and cc>=220 and cc<224) then grbp<="010";
	end if;
	if (ll=389 and cc>=225 and cc<247) then grbp<="010";
	end if;
	if (cc=13 and ll=390) then grbp<="010";
	end if;
	if (cc=15 and ll=390) then grbp<="010";
	end if;
	if (ll=390 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=390 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (ll=390 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (cc=100 and ll=390) then grbp<="010";
	end if;
	if (ll=390 and cc>=100 and cc<110) then grbp<="010";
	end if;
	if (ll=390 and cc>=112 and cc<154) then grbp<="010";
	end if;
	if (ll=390 and cc>=182 and cc<194) then grbp<="010";
	end if;
	if (ll=390 and cc>=203 and cc<208) then grbp<="010";
	end if;
	if (cc=220 and ll=390) then grbp<="010";
	end if;
	if (ll=390 and cc>=220 and cc<223) then grbp<="010";
	end if;
	if (ll=390 and cc>=225 and cc<247) then grbp<="010";
	end if;
	if (cc=13 and ll=391) then grbp<="010";
	end if;
	if (cc=15 and ll=391) then grbp<="010";
	end if;
	if (ll=391 and cc>=15 and cc<18) then grbp<="010";
	end if;
	if (ll=391 and cc>=30 and cc<36) then grbp<="010";
	end if;
	if (ll=391 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (cc=99 and ll=391) then grbp<="010";
	end if;
	if (ll=391 and cc>=99 and cc<110) then grbp<="010";
	end if;
	if (ll=391 and cc>=112 and cc<154) then grbp<="010";
	end if;
	if (ll=391 and cc>=182 and cc<195) then grbp<="010";
	end if;
	if (ll=391 and cc>=204 and cc<207) then grbp<="010";
	end if;
	if (ll=391 and cc>=219 and cc<223) then grbp<="010";
	end if;
	if (ll=391 and cc>=225 and cc<247) then grbp<="010";
	end if;
	if (cc=13 and ll=392) then grbp<="010";
	end if;
	if (cc=15 and ll=392) then grbp<="010";
	end if;
	if (ll=392 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=392 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=99 and ll=392) then grbp<="010";
	end if;
	if (ll=392 and cc>=99 and cc<109) then grbp<="010";
	end if;
	if (ll=392 and cc>=112 and cc<153) then grbp<="010";
	end if;
	if (ll=392 and cc>=183 and cc<195) then grbp<="010";
	end if;
	if (ll=392 and cc>=205 and cc<207) then grbp<="010";
	end if;
	if (ll=392 and cc>=219 and cc<222) then grbp<="010";
	end if;
	if (ll=392 and cc>=224 and cc<246) then grbp<="010";
	end if;
	if (cc=13 and ll=393) then grbp<="010";
	end if;
	if (cc=15 and ll=393) then grbp<="010";
	end if;
	if (ll=393 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=393 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (ll=393 and cc>=98 and cc<109) then grbp<="010";
	end if;
	if (ll=393 and cc>=111 and cc<152) then grbp<="010";
	end if;
	if (cc=183 and ll=393) then grbp<="010";
	end if;
	if (ll=393 and cc>=183 and cc<196) then grbp<="010";
	end if;
	if (cc=219 and ll=393) then grbp<="010";
	end if;
	if (ll=393 and cc>=219 and cc<222) then grbp<="010";
	end if;
	if (ll=393 and cc>=224 and cc<246) then grbp<="010";
	end if;
	if (ll=394 and cc>=1 and cc<3) then grbp<="010";
	end if;
	if (ll=394 and cc>=5 and cc<7) then grbp<="010";
	end if;
	if (cc=15 and ll=394) then grbp<="010";
	end if;
	if (ll=394 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=394 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=81 and ll=394) then grbp<="010";
	end if;
	if (cc=98 and ll=394) then grbp<="010";
	end if;
	if (ll=394 and cc>=98 and cc<108) then grbp<="010";
	end if;
	if (ll=394 and cc>=111 and cc<154) then grbp<="010";
	end if;
	if (ll=394 and cc>=183 and cc<197) then grbp<="010";
	end if;
	if (cc=211 and ll=394) then grbp<="010";
	end if;
	if (cc=218 and ll=394) then grbp<="010";
	end if;
	if (ll=394 and cc>=218 and cc<221) then grbp<="010";
	end if;
	if (ll=394 and cc>=224 and cc<246) then grbp<="010";
	end if;
	if (ll=395 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (cc=15 and ll=395) then grbp<="010";
	end if;
	if (ll=395 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=395 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=80 and ll=395) then grbp<="010";
	end if;
	if (ll=395 and cc>=80 and cc<82) then grbp<="010";
	end if;
	if (ll=395 and cc>=97 and cc<108) then grbp<="010";
	end if;
	if (ll=395 and cc>=111 and cc<153) then grbp<="010";
	end if;
	if (ll=395 and cc>=183 and cc<197) then grbp<="010";
	end if;
	if (cc=218 and ll=395) then grbp<="010";
	end if;
	if (ll=395 and cc>=218 and cc<220) then grbp<="010";
	end if;
	if (ll=395 and cc>=224 and cc<246) then grbp<="010";
	end if;
	if (ll=396 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (cc=15 and ll=396) then grbp<="010";
	end if;
	if (ll=396 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=396 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=97 and ll=396) then grbp<="010";
	end if;
	if (ll=396 and cc>=97 and cc<107) then grbp<="010";
	end if;
	if (ll=396 and cc>=110 and cc<154) then grbp<="010";
	end if;
	if (cc=183 and ll=396) then grbp<="010";
	end if;
	if (ll=396 and cc>=183 and cc<198) then grbp<="010";
	end if;
	if (cc=218 and ll=396) then grbp<="010";
	end if;
	if (cc=223 and ll=396) then grbp<="010";
	end if;
	if (ll=396 and cc>=223 and cc<246) then grbp<="010";
	end if;
	if (ll=397 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=397 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=397 and cc>=30 and cc<35) then grbp<="010";
	end if;
	if (ll=397 and cc>=97 and cc<107) then grbp<="010";
	end if;
	if (ll=397 and cc>=110 and cc<155) then grbp<="010";
	end if;
	if (cc=183 and ll=397) then grbp<="010";
	end if;
	if (ll=397 and cc>=183 and cc<198) then grbp<="010";
	end if;
	if (cc=217 and ll=397) then grbp<="010";
	end if;
	if (ll=397 and cc>=217 and cc<219) then grbp<="010";
	end if;
	if (ll=397 and cc>=223 and cc<247) then grbp<="010";
	end if;
	if (ll=398 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=398 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=398 and cc>=30 and cc<35) then grbp<="010";
	end if;
	if (cc=96 and ll=398) then grbp<="010";
	end if;
	if (ll=398 and cc>=96 and cc<106) then grbp<="010";
	end if;
	if (ll=398 and cc>=109 and cc<156) then grbp<="010";
	end if;
	if (ll=398 and cc>=184 and cc<199) then grbp<="010";
	end if;
	if (cc=217 and ll=398) then grbp<="010";
	end if;
	if (cc=223 and ll=398) then grbp<="010";
	end if;
	if (ll=398 and cc>=223 and cc<247) then grbp<="010";
	end if;
	if (ll=399 and cc>=0 and cc<7) then grbp<="010";
	end if;
	if (ll=399 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=399 and cc>=30 and cc<35) then grbp<="010";
	end if;
	if (ll=399 and cc>=76 and cc<78) then grbp<="010";
	end if;
	if (ll=399 and cc>=96 and cc<105) then grbp<="010";
	end if;
	if (ll=399 and cc>=109 and cc<156) then grbp<="010";
	end if;
	if (ll=399 and cc>=184 and cc<199) then grbp<="010";
	end if;
	if (cc=216 and ll=399) then grbp<="010";
	end if;
	if (ll=399 and cc>=216 and cc<218) then grbp<="010";
	end if;
	if (ll=399 and cc>=222 and cc<233) then grbp<="010";
	end if;
	if (ll=399 and cc>=234 and cc<247) then grbp<="010";
	end if;
	if (ll=400 and cc>=0 and cc<6) then grbp<="010";
	end if;
	if (ll=400 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=400 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (ll=400 and cc>=95 and cc<105) then grbp<="010";
	end if;
	if (ll=400 and cc>=108 and cc<156) then grbp<="010";
	end if;
	if (ll=400 and cc>=184 and cc<199) then grbp<="010";
	end if;
	if (cc=215 and ll=400) then grbp<="010";
	end if;
	if (ll=400 and cc>=215 and cc<217) then grbp<="010";
	end if;
	if (cc=225 and ll=400) then grbp<="010";
	end if;
	if (ll=400 and cc>=225 and cc<233) then grbp<="010";
	end if;
	if (ll=400 and cc>=234 and cc<246) then grbp<="010";
	end if;
	if (ll=401 and cc>=0 and cc<6) then grbp<="010";
	end if;
	if (ll=401 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=401 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=95 and ll=401) then grbp<="010";
	end if;
	if (ll=401 and cc>=95 and cc<104) then grbp<="010";
	end if;
	if (ll=401 and cc>=107 and cc<157) then grbp<="010";
	end if;
	if (ll=401 and cc>=184 and cc<201) then grbp<="010";
	end if;
	if (ll=401 and cc>=204 and cc<206) then grbp<="010";
	end if;
	if (ll=401 and cc>=214 and cc<217) then grbp<="010";
	end if;
	if (cc=225 and ll=401) then grbp<="010";
	end if;
	if (ll=401 and cc>=225 and cc<233) then grbp<="010";
	end if;
	if (ll=401 and cc>=234 and cc<246) then grbp<="010";
	end if;
	if (ll=402 and cc>=1 and cc<6) then grbp<="010";
	end if;
	if (ll=402 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=402 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=80 and ll=402) then grbp<="010";
	end if;
	if (cc=95 and ll=402) then grbp<="010";
	end if;
	if (ll=402 and cc>=95 and cc<103) then grbp<="010";
	end if;
	if (ll=402 and cc>=106 and cc<158) then grbp<="010";
	end if;
	if (ll=402 and cc>=184 and cc<206) then grbp<="010";
	end if;
	if (ll=402 and cc>=213 and cc<216) then grbp<="010";
	end if;
	if (ll=402 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=402 and cc>=225 and cc<233) then grbp<="010";
	end if;
	if (ll=402 and cc>=234 and cc<245) then grbp<="010";
	end if;
	if (ll=403 and cc>=1 and cc<6) then grbp<="010";
	end if;
	if (ll=403 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=403 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=95 and ll=403) then grbp<="010";
	end if;
	if (ll=403 and cc>=95 and cc<102) then grbp<="010";
	end if;
	if (ll=403 and cc>=105 and cc<131) then grbp<="010";
	end if;
	if (ll=403 and cc>=132 and cc<151) then grbp<="010";
	end if;
	if (cc=155 and ll=403) then grbp<="010";
	end if;
	if (ll=403 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (ll=403 and cc>=184 and cc<206) then grbp<="010";
	end if;
	if (ll=403 and cc>=213 and cc<216) then grbp<="010";
	end if;
	if (ll=403 and cc>=221 and cc<232) then grbp<="010";
	end if;
	if (ll=403 and cc>=234 and cc<245) then grbp<="010";
	end if;
	if (ll=404 and cc>=1 and cc<7) then grbp<="010";
	end if;
	if (ll=404 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=404 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (ll=404 and cc>=94 and cc<100) then grbp<="010";
	end if;
	if (ll=404 and cc>=104 and cc<131) then grbp<="010";
	end if;
	if (ll=404 and cc>=132 and cc<136) then grbp<="010";
	end if;
	if (cc=139 and ll=404) then grbp<="010";
	end if;
	if (ll=404 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (cc=155 and ll=404) then grbp<="010";
	end if;
	if (ll=404 and cc>=155 and cc<158) then grbp<="010";
	end if;
	if (ll=404 and cc>=185 and cc<201) then grbp<="010";
	end if;
	if (ll=404 and cc>=202 and cc<206) then grbp<="010";
	end if;
	if (cc=214 and ll=404) then grbp<="010";
	end if;
	if (cc=217 and ll=404) then grbp<="010";
	end if;
	if (ll=404 and cc>=217 and cc<221) then grbp<="010";
	end if;
	if (ll=404 and cc>=223 and cc<225) then grbp<="010";
	end if;
	if (ll=404 and cc>=228 and cc<232) then grbp<="010";
	end if;
	if (ll=404 and cc>=236 and cc<238) then grbp<="010";
	end if;
	if (ll=404 and cc>=241 and cc<243) then grbp<="010";
	end if;
	if (ll=405 and cc>=1 and cc<7) then grbp<="010";
	end if;
	if (ll=405 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=405 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=65 and ll=405) then grbp<="010";
	end if;
	if (cc=94 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=405 and cc>=103 and cc<131) then grbp<="010";
	end if;
	if (ll=405 and cc>=132 and cc<136) then grbp<="010";
	end if;
	if (cc=139 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=139 and cc<151) then grbp<="010";
	end if;
	if (cc=155 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=155 and cc<157) then grbp<="010";
	end if;
	if (ll=405 and cc>=185 and cc<199) then grbp<="010";
	end if;
	if (cc=202 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=202 and cc<206) then grbp<="010";
	end if;
	if (cc=219 and ll=405) then grbp<="010";
	end if;
	if (cc=221 and ll=405) then grbp<="010";
	end if;
	if (cc=223 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=223 and cc<225) then grbp<="010";
	end if;
	if (cc=228 and ll=405) then grbp<="010";
	end if;
	if (ll=405 and cc>=228 and cc<230) then grbp<="010";
	end if;
	if (cc=233 and ll=405) then grbp<="010";
	end if;
	if (cc=235 and ll=405) then grbp<="010";
	end if;
	if (cc=237 and ll=405) then grbp<="010";
	end if;
	if (cc=239 and ll=405) then grbp<="010";
	end if;
	if (cc=241 and ll=405) then grbp<="010";
	end if;
	if (cc=243 and ll=405) then grbp<="010";
	end if;
	if (cc=245 and ll=405) then grbp<="010";
	end if;
	if (cc=2 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=2 and cc<7) then grbp<="010";
	end if;
	if (ll=406 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=406 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (ll=406 and cc>=59 and cc<61) then grbp<="010";
	end if;
	if (cc=94 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=94 and cc<96) then grbp<="010";
	end if;
	if (ll=406 and cc>=102 and cc<131) then grbp<="010";
	end if;
	if (cc=139 and ll=406) then grbp<="010";
	end if;
	if (cc=143 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (cc=149 and ll=406) then grbp<="010";
	end if;
	if (cc=157 and ll=406) then grbp<="010";
	end if;
	if (cc=186 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=186 and cc<191) then grbp<="010";
	end if;
	if (ll=406 and cc>=192 and cc<195) then grbp<="010";
	end if;
	if (cc=200 and ll=406) then grbp<="010";
	end if;
	if (cc=202 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=202 and cc<205) then grbp<="010";
	end if;
	if (cc=214 and ll=406) then grbp<="010";
	end if;
	if (cc=216 and ll=406) then grbp<="010";
	end if;
	if (cc=219 and ll=406) then grbp<="010";
	end if;
	if (cc=222 and ll=406) then grbp<="010";
	end if;
	if (cc=226 and ll=406) then grbp<="010";
	end if;
	if (cc=228 and ll=406) then grbp<="010";
	end if;
	if (cc=231 and ll=406) then grbp<="010";
	end if;
	if (cc=234 and ll=406) then grbp<="010";
	end if;
	if (ll=406 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (ll=406 and cc>=237 and cc<240) then grbp<="010";
	end if;
	if (cc=244 and ll=406) then grbp<="010";
	end if;
	if (cc=2 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=2 and cc<7) then grbp<="010";
	end if;
	if (ll=407 and cc>=13 and cc<19) then grbp<="010";
	end if;
	if (ll=407 and cc>=30 and cc<34) then grbp<="010";
	end if;
	if (cc=100 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=100 and cc<131) then grbp<="010";
	end if;
	if (cc=143 and ll=407) then grbp<="010";
	end if;
	if (cc=147 and ll=407) then grbp<="010";
	end if;
	if (cc=149 and ll=407) then grbp<="010";
	end if;
	if (cc=151 and ll=407) then grbp<="010";
	end if;
	if (cc=153 and ll=407) then grbp<="010";
	end if;
	if (cc=187 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (cc=197 and ll=407) then grbp<="010";
	end if;
	if (cc=200 and ll=407) then grbp<="010";
	end if;
	if (cc=203 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (cc=210 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=407 and cc>=214 and cc<216) then grbp<="010";
	end if;
	if (cc=219 and ll=407) then grbp<="010";
	end if;
	if (cc=221 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=407 and cc>=227 and cc<230) then grbp<="010";
	end if;
	if (cc=234 and ll=407) then grbp<="010";
	end if;
	if (cc=236 and ll=407) then grbp<="010";
	end if;
	if (ll=407 and cc>=236 and cc<240) then grbp<="010";
	end if;
	if (cc=3 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=3 and cc<7) then grbp<="010";
	end if;
	if (ll=408 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (ll=408 and cc>=30 and cc<33) then grbp<="010";
	end if;
	if (ll=408 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (cc=79 and ll=408) then grbp<="010";
	end if;
	if (cc=99 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=99 and cc<131) then grbp<="010";
	end if;
	if (ll=408 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=408) then grbp<="010";
	end if;
	if (cc=139 and ll=408) then grbp<="010";
	end if;
	if (cc=141 and ll=408) then grbp<="010";
	end if;
	if (cc=143 and ll=408) then grbp<="010";
	end if;
	if (cc=145 and ll=408) then grbp<="010";
	end if;
	if (cc=147 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (cc=153 and ll=408) then grbp<="010";
	end if;
	if (cc=155 and ll=408) then grbp<="010";
	end if;
	if (cc=185 and ll=408) then grbp<="010";
	end if;
	if (cc=187 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (cc=193 and ll=408) then grbp<="010";
	end if;
	if (cc=195 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=195 and cc<197) then grbp<="010";
	end if;
	if (cc=200 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=200 and cc<202) then grbp<="010";
	end if;
	if (ll=408 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (cc=210 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=408 and cc>=214 and cc<216) then grbp<="010";
	end if;
	if (cc=219 and ll=408) then grbp<="010";
	end if;
	if (cc=221 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=408 and cc>=228 and cc<230) then grbp<="010";
	end if;
	if (cc=237 and ll=408) then grbp<="010";
	end if;
	if (ll=408 and cc>=237 and cc<239) then grbp<="010";
	end if;
	if (cc=4 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=4 and cc<7) then grbp<="010";
	end if;
	if (ll=409 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (ll=409 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=58 and ll=409) then grbp<="010";
	end if;
	if (cc=60 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (cc=97 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=97 and cc<131) then grbp<="010";
	end if;
	if (ll=409 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=409) then grbp<="010";
	end if;
	if (cc=139 and ll=409) then grbp<="010";
	end if;
	if (cc=141 and ll=409) then grbp<="010";
	end if;
	if (cc=143 and ll=409) then grbp<="010";
	end if;
	if (cc=147 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (cc=153 and ll=409) then grbp<="010";
	end if;
	if (cc=155 and ll=409) then grbp<="010";
	end if;
	if (cc=185 and ll=409) then grbp<="010";
	end if;
	if (cc=187 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (cc=193 and ll=409) then grbp<="010";
	end if;
	if (cc=198 and ll=409) then grbp<="010";
	end if;
	if (cc=201 and ll=409) then grbp<="010";
	end if;
	if (cc=203 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (cc=208 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (ll=409 and cc>=214 and cc<218) then grbp<="010";
	end if;
	if (cc=221 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=409 and cc>=225 and cc<227) then grbp<="010";
	end if;
	if (cc=231 and ll=409) then grbp<="010";
	end if;
	if (cc=234 and ll=409) then grbp<="010";
	end if;
	if (ll=409 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (ll=409 and cc>=237 and cc<240) then grbp<="010";
	end if;
	if (cc=4 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=4 and cc<8) then grbp<="010";
	end if;
	if (ll=410 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (cc=54 and ll=410) then grbp<="010";
	end if;
	if (cc=58 and ll=410) then grbp<="010";
	end if;
	if (cc=66 and ll=410) then grbp<="010";
	end if;
	if (cc=80 and ll=410) then grbp<="010";
	end if;
	if (cc=95 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=95 and cc<131) then grbp<="010";
	end if;
	if (ll=410 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=410) then grbp<="010";
	end if;
	if (cc=139 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=410 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (ll=410 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (cc=153 and ll=410) then grbp<="010";
	end if;
	if (cc=155 and ll=410) then grbp<="010";
	end if;
	if (cc=187 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=187 and cc<190) then grbp<="010";
	end if;
	if (cc=193 and ll=410) then grbp<="010";
	end if;
	if (cc=195 and ll=410) then grbp<="010";
	end if;
	if (cc=197 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=197 and cc<199) then grbp<="010";
	end if;
	if (cc=203 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (cc=208 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=208 and cc<213) then grbp<="010";
	end if;
	if (cc=219 and ll=410) then grbp<="010";
	end if;
	if (cc=221 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=410 and cc>=225 and cc<227) then grbp<="010";
	end if;
	if (cc=234 and ll=410) then grbp<="010";
	end if;
	if (ll=410 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (ll=410 and cc>=238 and cc<240) then grbp<="010";
	end if;
	if (ll=411 and cc>=5 and cc<8) then grbp<="010";
	end if;
	if (ll=411 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (ll=411 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=65 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=65 and cc<68) then grbp<="010";
	end if;
	if (ll=411 and cc>=93 and cc<131) then grbp<="010";
	end if;
	if (ll=411 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=411) then grbp<="010";
	end if;
	if (cc=139 and ll=411) then grbp<="010";
	end if;
	if (cc=141 and ll=411) then grbp<="010";
	end if;
	if (cc=143 and ll=411) then grbp<="010";
	end if;
	if (cc=145 and ll=411) then grbp<="010";
	end if;
	if (cc=147 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (cc=155 and ll=411) then grbp<="010";
	end if;
	if (cc=187 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=187 and cc<192) then grbp<="010";
	end if;
	if (cc=195 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=195 and cc<197) then grbp<="010";
	end if;
	if (cc=203 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=203 and cc<205) then grbp<="010";
	end if;
	if (cc=208 and ll=411) then grbp<="010";
	end if;
	if (cc=210 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=411 and cc>=214 and cc<218) then grbp<="010";
	end if;
	if (cc=221 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=221 and cc<223) then grbp<="010";
	end if;
	if (ll=411 and cc>=225 and cc<227) then grbp<="010";
	end if;
	if (cc=234 and ll=411) then grbp<="010";
	end if;
	if (ll=411 and cc>=234 and cc<236) then grbp<="010";
	end if;
	if (cc=241 and ll=411) then grbp<="010";
	end if;
	if (cc=244 and ll=411) then grbp<="010";
	end if;
	if (cc=6 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=6 and cc<8) then grbp<="010";
	end if;
	if (ll=412 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (ll=412 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=72 and ll=412) then grbp<="010";
	end if;
	if (cc=80 and ll=412) then grbp<="010";
	end if;
	if (cc=92 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=92 and cc<131) then grbp<="010";
	end if;
	if (ll=412 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=412) then grbp<="010";
	end if;
	if (cc=143 and ll=412) then grbp<="010";
	end if;
	if (cc=147 and ll=412) then grbp<="010";
	end if;
	if (cc=150 and ll=412) then grbp<="010";
	end if;
	if (cc=152 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=152 and cc<154) then grbp<="010";
	end if;
	if (cc=187 and ll=412) then grbp<="010";
	end if;
	if (cc=189 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=189 and cc<192) then grbp<="010";
	end if;
	if (cc=197 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=197 and cc<199) then grbp<="010";
	end if;
	if (ll=412 and cc>=201 and cc<203) then grbp<="010";
	end if;
	if (cc=210 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=210 and cc<213) then grbp<="010";
	end if;
	if (ll=412 and cc>=214 and cc<218) then grbp<="010";
	end if;
	if (cc=223 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=223 and cc<225) then grbp<="010";
	end if;
	if (cc=232 and ll=412) then grbp<="010";
	end if;
	if (ll=412 and cc>=232 and cc<234) then grbp<="010";
	end if;
	if (cc=242 and ll=412) then grbp<="010";
	end if;
	if (cc=7 and ll=413) then grbp<="010";
	end if;
	if (cc=14 and ll=413) then grbp<="010";
	end if;
	if (ll=413 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (ll=413 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=62 and ll=413) then grbp<="010";
	end if;
	if (cc=66 and ll=413) then grbp<="010";
	end if;
	if (cc=72 and ll=413) then grbp<="010";
	end if;
	if (cc=92 and ll=413) then grbp<="010";
	end if;
	if (ll=413 and cc>=92 and cc<131) then grbp<="010";
	end if;
	if (ll=413 and cc>=132 and cc<134) then grbp<="010";
	end if;
	if (cc=137 and ll=413) then grbp<="010";
	end if;
	if (cc=139 and ll=413) then grbp<="010";
	end if;
	if (cc=142 and ll=413) then grbp<="010";
	end if;
	if (ll=413 and cc>=142 and cc<144) then grbp<="010";
	end if;
	if (cc=149 and ll=413) then grbp<="010";
	end if;
	if (ll=413 and cc>=149 and cc<151) then grbp<="010";
	end if;
	if (ll=413 and cc>=152 and cc<154) then grbp<="010";
	end if;
	if (cc=159 and ll=413) then grbp<="010";
	end if;
	if (ll=413 and cc>=159 and cc<161) then grbp<="010";
	end if;
	if (ll=413 and cc>=186 and cc<195) then grbp<="010";
	end if;
	if (ll=413 and cc>=197 and cc<199) then grbp<="010";
	end if;
	if (ll=413 and cc>=200 and cc<208) then grbp<="010";
	end if;
	if (ll=413 and cc>=209 and cc<221) then grbp<="010";
	end if;
	if (ll=413 and cc>=222 and cc<231) then grbp<="010";
	end if;
	if (ll=413 and cc>=232 and cc<234) then grbp<="010";
	end if;
	if (ll=413 and cc>=236 and cc<238) then grbp<="010";
	end if;
	if (ll=413 and cc>=240 and cc<242) then grbp<="010";
	end if;
	if (ll=413 and cc>=243 and cc<245) then grbp<="010";
	end if;
	if (cc=14 and ll=414) then grbp<="010";
	end if;
	if (ll=414 and cc>=14 and cc<19) then grbp<="010";
	end if;
	if (cc=72 and ll=414) then grbp<="010";
	end if;
	if (cc=91 and ll=414) then grbp<="010";
	end if;
	if (ll=414 and cc>=91 and cc<140) then grbp<="010";
	end if;
	if (ll=414 and cc>=141 and cc<160) then grbp<="010";
	end if;
	if (cc=188 and ll=414) then grbp<="010";
	end if;
	if (ll=414 and cc>=188 and cc<225) then grbp<="010";
	end if;
	if (cc=232 and ll=414) then grbp<="010";
	end if;
	if (ll=414 and cc>=232 and cc<242) then grbp<="010";
	end if;
	if (cc=15 and ll=415) then grbp<="010";
	end if;
	if (ll=415 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=415 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=91 and ll=415) then grbp<="010";
	end if;
	if (ll=415 and cc>=91 and cc<140) then grbp<="010";
	end if;
	if (ll=415 and cc>=141 and cc<160) then grbp<="010";
	end if;
	if (cc=188 and ll=415) then grbp<="010";
	end if;
	if (ll=415 and cc>=188 and cc<225) then grbp<="010";
	end if;
	if (cc=231 and ll=415) then grbp<="010";
	end if;
	if (ll=415 and cc>=231 and cc<242) then grbp<="010";
	end if;
	if (cc=15 and ll=416) then grbp<="010";
	end if;
	if (ll=416 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=416 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=73 and ll=416) then grbp<="010";
	end if;
	if (cc=78 and ll=416) then grbp<="010";
	end if;
	if (cc=90 and ll=416) then grbp<="010";
	end if;
	if (ll=416 and cc>=90 and cc<160) then grbp<="010";
	end if;
	if (ll=416 and cc>=188 and cc<225) then grbp<="010";
	end if;
	if (ll=416 and cc>=229 and cc<241) then grbp<="010";
	end if;
	if (cc=7 and ll=417) then grbp<="010";
	end if;
	if (cc=15 and ll=417) then grbp<="010";
	end if;
	if (ll=417 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=417 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=79 and ll=417) then grbp<="010";
	end if;
	if (cc=89 and ll=417) then grbp<="010";
	end if;
	if (ll=417 and cc>=89 and cc<160) then grbp<="010";
	end if;
	if (ll=417 and cc>=188 and cc<225) then grbp<="010";
	end if;
	if (ll=417 and cc>=230 and cc<240) then grbp<="010";
	end if;
	if (cc=7 and ll=418) then grbp<="010";
	end if;
	if (cc=15 and ll=418) then grbp<="010";
	end if;
	if (ll=418 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=418 and cc>=30 and cc<32) then grbp<="010";
	end if;
	if (cc=89 and ll=418) then grbp<="010";
	end if;
	if (ll=418 and cc>=89 and cc<160) then grbp<="010";
	end if;
	if (ll=418 and cc>=189 and cc<225) then grbp<="010";
	end if;
	if (ll=418 and cc>=226 and cc<240) then grbp<="010";
	end if;
	if (cc=7 and ll=419) then grbp<="010";
	end if;
	if (cc=15 and ll=419) then grbp<="010";
	end if;
	if (ll=419 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=419 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=75 and ll=419) then grbp<="010";
	end if;
	if (cc=88 and ll=419) then grbp<="010";
	end if;
	if (ll=419 and cc>=88 and cc<156) then grbp<="010";
	end if;
	if (ll=419 and cc>=157 and cc<160) then grbp<="010";
	end if;
	if (cc=189 and ll=419) then grbp<="010";
	end if;
	if (ll=419 and cc>=189 and cc<227) then grbp<="010";
	end if;
	if (ll=419 and cc>=228 and cc<239) then grbp<="010";
	end if;
	if (ll=419 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=420) then grbp<="010";
	end if;
	if (cc=15 and ll=420) then grbp<="010";
	end if;
	if (ll=420 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=420 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=58 and ll=420) then grbp<="010";
	end if;
	if (cc=64 and ll=420) then grbp<="010";
	end if;
	if (cc=68 and ll=420) then grbp<="010";
	end if;
	if (cc=73 and ll=420) then grbp<="010";
	end if;
	if (cc=88 and ll=420) then grbp<="010";
	end if;
	if (ll=420 and cc>=88 and cc<158) then grbp<="010";
	end if;
	if (cc=187 and ll=420) then grbp<="010";
	end if;
	if (cc=189 and ll=420) then grbp<="010";
	end if;
	if (ll=420 and cc>=189 and cc<239) then grbp<="010";
	end if;
	if (ll=420 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=421) then grbp<="010";
	end if;
	if (cc=15 and ll=421) then grbp<="010";
	end if;
	if (ll=421 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=421 and cc>=29 and cc<32) then grbp<="010";
	end if;
	if (cc=58 and ll=421) then grbp<="010";
	end if;
	if (cc=68 and ll=421) then grbp<="010";
	end if;
	if (cc=79 and ll=421) then grbp<="010";
	end if;
	if (cc=87 and ll=421) then grbp<="010";
	end if;
	if (ll=421 and cc>=87 and cc<160) then grbp<="010";
	end if;
	if (cc=189 and ll=421) then grbp<="010";
	end if;
	if (ll=421 and cc>=189 and cc<221) then grbp<="010";
	end if;
	if (ll=421 and cc>=223 and cc<239) then grbp<="010";
	end if;
	if (ll=421 and cc>=248 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=422) then grbp<="010";
	end if;
	if (cc=15 and ll=422) then grbp<="010";
	end if;
	if (ll=422 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=422 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=61 and ll=422) then grbp<="010";
	end if;
	if (cc=83 and ll=422) then grbp<="010";
	end if;
	if (cc=87 and ll=422) then grbp<="010";
	end if;
	if (ll=422 and cc>=87 and cc<157) then grbp<="010";
	end if;
	if (cc=187 and ll=422) then grbp<="010";
	end if;
	if (ll=422 and cc>=187 and cc<220) then grbp<="010";
	end if;
	if (ll=422 and cc>=221 and cc<238) then grbp<="010";
	end if;
	if (ll=422 and cc>=247 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=423) then grbp<="010";
	end if;
	if (cc=15 and ll=423) then grbp<="010";
	end if;
	if (ll=423 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=423 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=86 and ll=423) then grbp<="010";
	end if;
	if (ll=423 and cc>=86 and cc<157) then grbp<="010";
	end if;
	if (cc=188 and ll=423) then grbp<="010";
	end if;
	if (ll=423 and cc>=188 and cc<219) then grbp<="010";
	end if;
	if (ll=423 and cc>=221 and cc<237) then grbp<="010";
	end if;
	if (ll=423 and cc>=247 and cc<251) then grbp<="010";
	end if;
	if (cc=7 and ll=424) then grbp<="010";
	end if;
	if (cc=15 and ll=424) then grbp<="010";
	end if;
	if (ll=424 and cc>=15 and cc<19) then grbp<="010";
	end if;
	if (ll=424 and cc>=29 and cc<31) then grbp<="010";
	end if;
	if (cc=86 and ll=424) then grbp<="010";
	end if;
	if (ll=424 and cc>=86 and cc<157) then grbp<="010";
	end if;
	if (cc=189 and ll=424) then grbp<="010";
	end if;
	if (ll=424 and cc>=189 and cc<219) then grbp<="010";
	end if;
	if (ll=424 and cc>=221 and cc<237) then grbp<="010";
	end if;
	if (ll=424 and cc>=247 and cc<251) then grbp<="010";
	end if;


	if (cc=0 and ll=0) then grbp<="110";
	end if;
	if (cc=2 and ll=0) then grbp<="110";
	end if;
	if (ll=0 and cc>=2 and cc<13) then grbp<="110";
	end if;
	if (ll=0 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=0 and cc>=164 and cc<169) then grbp<="110";
	end if;
	if (ll=0 and cc>=172 and cc<179) then grbp<="110";
	end if;
	if (cc=182 and ll=0) then grbp<="110";
	end if;
	if (cc=186 and ll=0) then grbp<="110";
	end if;
	if (ll=0 and cc>=186 and cc<198) then grbp<="110";
	end if;
	if (cc=249 and ll=0) then grbp<="110";
	end if;
	if (cc=0 and ll=1) then grbp<="110";
	end if;
	if (cc=2 and ll=1) then grbp<="110";
	end if;
	if (ll=1 and cc>=2 and cc<13) then grbp<="110";
	end if;
	if (ll=1 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=1 and cc>=164 and cc<169) then grbp<="110";
	end if;
	if (ll=1 and cc>=172 and cc<179) then grbp<="110";
	end if;
	if (cc=182 and ll=1) then grbp<="110";
	end if;
	if (cc=186 and ll=1) then grbp<="110";
	end if;
	if (ll=1 and cc>=186 and cc<198) then grbp<="110";
	end if;
	if (cc=249 and ll=1) then grbp<="110";
	end if;
	if (cc=0 and ll=2) then grbp<="110";
	end if;
	if (cc=2 and ll=2) then grbp<="110";
	end if;
	if (ll=2 and cc>=2 and cc<13) then grbp<="110";
	end if;
	if (ll=2 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=2 and cc>=164 and cc<169) then grbp<="110";
	end if;
	if (ll=2 and cc>=172 and cc<179) then grbp<="110";
	end if;
	if (cc=182 and ll=2) then grbp<="110";
	end if;
	if (cc=186 and ll=2) then grbp<="110";
	end if;
	if (ll=2 and cc>=186 and cc<198) then grbp<="110";
	end if;
	if (cc=249 and ll=2) then grbp<="110";
	end if;
	if (cc=0 and ll=3) then grbp<="110";
	end if;
	if (cc=2 and ll=3) then grbp<="110";
	end if;
	if (ll=3 and cc>=2 and cc<13) then grbp<="110";
	end if;
	if (ll=3 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=3 and cc>=164 and cc<169) then grbp<="110";
	end if;
	if (ll=3 and cc>=172 and cc<179) then grbp<="110";
	end if;
	if (cc=182 and ll=3) then grbp<="110";
	end if;
	if (cc=186 and ll=3) then grbp<="110";
	end if;
	if (ll=3 and cc>=186 and cc<198) then grbp<="110";
	end if;
	if (cc=249 and ll=3) then grbp<="110";
	end if;
	if (cc=0 and ll=4) then grbp<="110";
	end if;
	if (ll=4 and cc>=0 and cc<6) then grbp<="110";
	end if;
	if (ll=4 and cc>=7 and cc<10) then grbp<="110";
	end if;
	if (ll=4 and cc>=12 and cc<14) then grbp<="110";
	end if;
	if (cc=17 and ll=4) then grbp<="110";
	end if;
	if (ll=4 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=4 and cc>=164 and cc<168) then grbp<="110";
	end if;
	if (cc=173 and ll=4) then grbp<="110";
	end if;
	if (cc=175 and ll=4) then grbp<="110";
	end if;
	if (ll=4 and cc>=175 and cc<180) then grbp<="110";
	end if;
	if (ll=4 and cc>=186 and cc<189) then grbp<="110";
	end if;
	if (ll=4 and cc>=190 and cc<196) then grbp<="110";
	end if;
	if (ll=4 and cc>=197 and cc<199) then grbp<="110";
	end if;
	if (ll=5 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (cc=12 and ll=5) then grbp<="110";
	end if;
	if (ll=5 and cc>=12 and cc<14) then grbp<="110";
	end if;
	if (ll=5 and cc>=15 and cc<27) then grbp<="110";
	end if;
	if (ll=5 and cc>=164 and cc<169) then grbp<="110";
	end if;
	if (ll=5 and cc>=173 and cc<175) then grbp<="110";
	end if;
	if (ll=5 and cc>=176 and cc<179) then grbp<="110";
	end if;
	if (ll=5 and cc>=183 and cc<186) then grbp<="110";
	end if;
	if (ll=5 and cc>=188 and cc<196) then grbp<="110";
	end if;
	if (ll=5 and cc>=197 and cc<199) then grbp<="110";
	end if;
	if (cc=0 and ll=6) then grbp<="110";
	end if;
	if (ll=6 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=6 and cc>=9 and cc<11) then grbp<="110";
	end if;
	if (cc=16 and ll=6) then grbp<="110";
	end if;
	if (ll=6 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (ll=6 and cc>=163 and cc<170) then grbp<="110";
	end if;
	if (ll=6 and cc>=173 and cc<176) then grbp<="110";
	end if;
	if (ll=6 and cc>=178 and cc<183) then grbp<="110";
	end if;
	if (cc=186 and ll=6) then grbp<="110";
	end if;
	if (cc=188 and ll=6) then grbp<="110";
	end if;
	if (ll=6 and cc>=188 and cc<197) then grbp<="110";
	end if;
	if (cc=207 and ll=6) then grbp<="110";
	end if;
	if (cc=0 and ll=7) then grbp<="110";
	end if;
	if (ll=7 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=7 and cc>=8 and cc<11) then grbp<="110";
	end if;
	if (ll=7 and cc>=12 and cc<14) then grbp<="110";
	end if;
	if (cc=17 and ll=7) then grbp<="110";
	end if;
	if (ll=7 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=7 and cc>=165 and cc<172) then grbp<="110";
	end if;
	if (ll=7 and cc>=173 and cc<183) then grbp<="110";
	end if;
	if (ll=7 and cc>=184 and cc<186) then grbp<="110";
	end if;
	if (ll=7 and cc>=187 and cc<197) then grbp<="110";
	end if;
	if (ll=7 and cc>=198 and cc<200) then grbp<="110";
	end if;
	if (cc=0 and ll=8) then grbp<="110";
	end if;
	if (ll=8 and cc>=0 and cc<3) then grbp<="110";
	end if;
	if (ll=8 and cc>=4 and cc<7) then grbp<="110";
	end if;
	if (ll=8 and cc>=8 and cc<11) then grbp<="110";
	end if;
	if (ll=8 and cc>=13 and cc<16) then grbp<="110";
	end if;
	if (ll=8 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=8 and cc>=165 and cc<170) then grbp<="110";
	end if;
	if (cc=173 and ll=8) then grbp<="110";
	end if;
	if (ll=8 and cc>=173 and cc<187) then grbp<="110";
	end if;
	if (cc=191 and ll=8) then grbp<="110";
	end if;
	if (ll=8 and cc>=191 and cc<194) then grbp<="110";
	end if;
	if (ll=8 and cc>=195 and cc<197) then grbp<="110";
	end if;
	if (ll=8 and cc>=198 and cc<200) then grbp<="110";
	end if;
	if (cc=0 and ll=9) then grbp<="110";
	end if;
	if (ll=9 and cc>=0 and cc<3) then grbp<="110";
	end if;
	if (ll=9 and cc>=4 and cc<9) then grbp<="110";
	end if;
	if (cc=13 and ll=9) then grbp<="110";
	end if;
	if (cc=16 and ll=9) then grbp<="110";
	end if;
	if (ll=9 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (ll=9 and cc>=166 and cc<187) then grbp<="110";
	end if;
	if (cc=192 and ll=9) then grbp<="110";
	end if;
	if (ll=9 and cc>=192 and cc<195) then grbp<="110";
	end if;
	if (cc=199 and ll=9) then grbp<="110";
	end if;
	if (cc=208 and ll=9) then grbp<="110";
	end if;
	if (cc=0 and ll=10) then grbp<="110";
	end if;
	if (ll=10 and cc>=0 and cc<6) then grbp<="110";
	end if;
	if (ll=10 and cc>=7 and cc<13) then grbp<="110";
	end if;
	if (ll=10 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=10 and cc>=166 and cc<188) then grbp<="110";
	end if;
	if (ll=10 and cc>=189 and cc<191) then grbp<="110";
	end if;
	if (ll=10 and cc>=193 and cc<197) then grbp<="110";
	end if;
	if (ll=10 and cc>=199 and cc<201) then grbp<="110";
	end if;
	if (ll=11 and cc>=0 and cc<9) then grbp<="110";
	end if;
	if (ll=11 and cc>=10 and cc<27) then grbp<="110";
	end if;
	if (ll=11 and cc>=166 and cc<187) then grbp<="110";
	end if;
	if (cc=190 and ll=11) then grbp<="110";
	end if;
	if (cc=193 and ll=11) then grbp<="110";
	end if;
	if (ll=11 and cc>=193 and cc<196) then grbp<="110";
	end if;
	if (cc=209 and ll=11) then grbp<="110";
	end if;
	if (cc=0 and ll=12) then grbp<="110";
	end if;
	if (ll=12 and cc>=0 and cc<11) then grbp<="110";
	end if;
	if (ll=12 and cc>=12 and cc<27) then grbp<="110";
	end if;
	if (ll=12 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (ll=12 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (cc=196 and ll=12) then grbp<="110";
	end if;
	if (ll=12 and cc>=196 and cc<198) then grbp<="110";
	end if;
	if (ll=12 and cc>=200 and cc<202) then grbp<="110";
	end if;
	if (ll=13 and cc>=0 and cc<12) then grbp<="110";
	end if;
	if (ll=13 and cc>=13 and cc<27) then grbp<="110";
	end if;
	if (ll=13 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (ll=13 and cc>=189 and cc<191) then grbp<="110";
	end if;
	if (cc=194 and ll=13) then grbp<="110";
	end if;
	if (cc=200 and ll=13) then grbp<="110";
	end if;
	if (cc=210 and ll=13) then grbp<="110";
	end if;
	if (cc=0 and ll=14) then grbp<="110";
	end if;
	if (ll=14 and cc>=0 and cc<3) then grbp<="110";
	end if;
	if (ll=14 and cc>=4 and cc<8) then grbp<="110";
	end if;
	if (cc=11 and ll=14) then grbp<="110";
	end if;
	if (cc=14 and ll=14) then grbp<="110";
	end if;
	if (ll=14 and cc>=14 and cc<27) then grbp<="110";
	end if;
	if (ll=14 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (cc=189 and ll=14) then grbp<="110";
	end if;
	if (ll=14 and cc>=189 and cc<191) then grbp<="110";
	end if;
	if (cc=194 and ll=14) then grbp<="110";
	end if;
	if (cc=201 and ll=14) then grbp<="110";
	end if;
	if (cc=210 and ll=14) then grbp<="110";
	end if;
	if (cc=0 and ll=15) then grbp<="110";
	end if;
	if (ll=15 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (ll=15 and cc>=11 and cc<26) then grbp<="110";
	end if;
	if (ll=15 and cc>=166 and cc<187) then grbp<="110";
	end if;
	if (ll=15 and cc>=188 and cc<190) then grbp<="110";
	end if;
	if (cc=193 and ll=15) then grbp<="110";
	end if;
	if (cc=196 and ll=15) then grbp<="110";
	end if;
	if (cc=201 and ll=15) then grbp<="110";
	end if;
	if (cc=210 and ll=15) then grbp<="110";
	end if;
	if (cc=0 and ll=16) then grbp<="110";
	end if;
	if (ll=16 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (cc=13 and ll=16) then grbp<="110";
	end if;
	if (ll=16 and cc>=13 and cc<27) then grbp<="110";
	end if;
	if (ll=16 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (ll=16 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (cc=195 and ll=16) then grbp<="110";
	end if;
	if (cc=201 and ll=16) then grbp<="110";
	end if;
	if (ll=16 and cc>=201 and cc<203) then grbp<="110";
	end if;
	if (cc=0 and ll=17) then grbp<="110";
	end if;
	if (ll=17 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (cc=13 and ll=17) then grbp<="110";
	end if;
	if (ll=17 and cc>=13 and cc<27) then grbp<="110";
	end if;
	if (ll=17 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (ll=17 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (cc=202 and ll=17) then grbp<="110";
	end if;
	if (cc=211 and ll=17) then grbp<="110";
	end if;
	if (cc=0 and ll=18) then grbp<="110";
	end if;
	if (ll=18 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=18 and cc>=3 and cc<26) then grbp<="110";
	end if;
	if (ll=18 and cc>=167 and cc<183) then grbp<="110";
	end if;
	if (ll=18 and cc>=184 and cc<188) then grbp<="110";
	end if;
	if (cc=202 and ll=18) then grbp<="110";
	end if;
	if (cc=211 and ll=18) then grbp<="110";
	end if;
	if (cc=0 and ll=19) then grbp<="110";
	end if;
	if (ll=19 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=19 and cc>=3 and cc<10) then grbp<="110";
	end if;
	if (ll=19 and cc>=11 and cc<27) then grbp<="110";
	end if;
	if (ll=19 and cc>=167 and cc<184) then grbp<="110";
	end if;
	if (ll=19 and cc>=185 and cc<190) then grbp<="110";
	end if;
	if (cc=193 and ll=19) then grbp<="110";
	end if;
	if (ll=19 and cc>=193 and cc<195) then grbp<="110";
	end if;
	if (ll=19 and cc>=202 and cc<204) then grbp<="110";
	end if;
	if (cc=0 and ll=20) then grbp<="110";
	end if;
	if (cc=3 and ll=20) then grbp<="110";
	end if;
	if (ll=20 and cc>=3 and cc<26) then grbp<="110";
	end if;
	if (ll=20 and cc>=167 and cc<187) then grbp<="110";
	end if;
	if (ll=20 and cc>=188 and cc<190) then grbp<="110";
	end if;
	if (cc=203 and ll=20) then grbp<="110";
	end if;
	if (cc=212 and ll=20) then grbp<="110";
	end if;
	if (cc=0 and ll=21) then grbp<="110";
	end if;
	if (cc=2 and ll=21) then grbp<="110";
	end if;
	if (ll=21 and cc>=2 and cc<26) then grbp<="110";
	end if;
	if (ll=21 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (cc=193 and ll=21) then grbp<="110";
	end if;
	if (cc=203 and ll=21) then grbp<="110";
	end if;
	if (cc=0 and ll=22) then grbp<="110";
	end if;
	if (ll=22 and cc>=0 and cc<26) then grbp<="110";
	end if;
	if (ll=22 and cc>=167 and cc<186) then grbp<="110";
	end if;
	if (ll=22 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (ll=22 and cc>=192 and cc<195) then grbp<="110";
	end if;
	if (cc=203 and ll=22) then grbp<="110";
	end if;
	if (ll=22 and cc>=203 and cc<205) then grbp<="110";
	end if;
	if (cc=0 and ll=23) then grbp<="110";
	end if;
	if (ll=23 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=23 and cc>=167 and cc<191) then grbp<="110";
	end if;
	if (ll=23 and cc>=192 and cc<194) then grbp<="110";
	end if;
	if (cc=204 and ll=23) then grbp<="110";
	end if;
	if (cc=213 and ll=23) then grbp<="110";
	end if;
	if (cc=0 and ll=24) then grbp<="110";
	end if;
	if (ll=24 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=24 and cc>=168 and cc<187) then grbp<="110";
	end if;
	if (cc=190 and ll=24) then grbp<="110";
	end if;
	if (ll=24 and cc>=190 and cc<195) then grbp<="110";
	end if;
	if (ll=24 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (cc=0 and ll=25) then grbp<="110";
	end if;
	if (ll=25 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=25 and cc>=168 and cc<190) then grbp<="110";
	end if;
	if (ll=25 and cc>=191 and cc<194) then grbp<="110";
	end if;
	if (cc=204 and ll=25) then grbp<="110";
	end if;
	if (ll=25 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (cc=0 and ll=26) then grbp<="110";
	end if;
	if (ll=26 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=26 and cc>=168 and cc<198) then grbp<="110";
	end if;
	if (ll=26 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (ll=27 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=27 and cc>=169 and cc<187) then grbp<="110";
	end if;
	if (ll=27 and cc>=188 and cc<198) then grbp<="110";
	end if;
	if (ll=27 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (cc=0 and ll=28) then grbp<="110";
	end if;
	if (ll=28 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=28 and cc>=169 and cc<197) then grbp<="110";
	end if;
	if (cc=215 and ll=28) then grbp<="110";
	end if;
	if (cc=0 and ll=29) then grbp<="110";
	end if;
	if (ll=29 and cc>=0 and cc<26) then grbp<="110";
	end if;
	if (ll=29 and cc>=170 and cc<181) then grbp<="110";
	end if;
	if (ll=29 and cc>=182 and cc<191) then grbp<="110";
	end if;
	if (ll=29 and cc>=192 and cc<197) then grbp<="110";
	end if;
	if (cc=0 and ll=30) then grbp<="110";
	end if;
	if (ll=30 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=30 and cc>=170 and cc<183) then grbp<="110";
	end if;
	if (ll=30 and cc>=184 and cc<186) then grbp<="110";
	end if;
	if (ll=30 and cc>=187 and cc<191) then grbp<="110";
	end if;
	if (ll=30 and cc>=192 and cc<194) then grbp<="110";
	end if;
	if (ll=30 and cc>=195 and cc<197) then grbp<="110";
	end if;
	if (cc=216 and ll=30) then grbp<="110";
	end if;
	if (cc=0 and ll=31) then grbp<="110";
	end if;
	if (ll=31 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=31 and cc>=171 and cc<186) then grbp<="110";
	end if;
	if (ll=31 and cc>=187 and cc<194) then grbp<="110";
	end if;
	if (cc=207 and ll=31) then grbp<="110";
	end if;
	if (cc=216 and ll=31) then grbp<="110";
	end if;
	if (cc=0 and ll=32) then grbp<="110";
	end if;
	if (ll=32 and cc>=0 and cc<26) then grbp<="110";
	end if;
	if (ll=32 and cc>=172 and cc<186) then grbp<="110";
	end if;
	if (ll=32 and cc>=188 and cc<194) then grbp<="110";
	end if;
	if (cc=216 and ll=32) then grbp<="110";
	end if;
	if (cc=0 and ll=33) then grbp<="110";
	end if;
	if (ll=33 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (cc=173 and ll=33) then grbp<="110";
	end if;
	if (ll=33 and cc>=173 and cc<181) then grbp<="110";
	end if;
	if (cc=184 and ll=33) then grbp<="110";
	end if;
	if (ll=33 and cc>=184 and cc<186) then grbp<="110";
	end if;
	if (ll=33 and cc>=188 and cc<195) then grbp<="110";
	end if;
	if (cc=217 and ll=33) then grbp<="110";
	end if;
	if (cc=0 and ll=34) then grbp<="110";
	end if;
	if (ll=34 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (cc=173 and ll=34) then grbp<="110";
	end if;
	if (ll=34 and cc>=173 and cc<186) then grbp<="110";
	end if;
	if (ll=34 and cc>=188 and cc<195) then grbp<="110";
	end if;
	if (cc=217 and ll=34) then grbp<="110";
	end if;
	if (cc=0 and ll=35) then grbp<="110";
	end if;
	if (ll=35 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=35 and cc>=174 and cc<180) then grbp<="110";
	end if;
	if (ll=35 and cc>=181 and cc<183) then grbp<="110";
	end if;
	if (ll=35 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (ll=35 and cc>=191 and cc<194) then grbp<="110";
	end if;
	if (cc=217 and ll=35) then grbp<="110";
	end if;
	if (cc=0 and ll=36) then grbp<="110";
	end if;
	if (ll=36 and cc>=0 and cc<27) then grbp<="110";
	end if;
	if (ll=36 and cc>=175 and cc<179) then grbp<="110";
	end if;
	if (cc=183 and ll=36) then grbp<="110";
	end if;
	if (ll=36 and cc>=183 and cc<185) then grbp<="110";
	end if;
	if (ll=36 and cc>=186 and cc<189) then grbp<="110";
	end if;
	if (ll=36 and cc>=191 and cc<193) then grbp<="110";
	end if;
	if (cc=218 and ll=36) then grbp<="110";
	end if;
	if (cc=0 and ll=37) then grbp<="110";
	end if;
	if (ll=37 and cc>=0 and cc<12) then grbp<="110";
	end if;
	if (ll=37 and cc>=13 and cc<27) then grbp<="110";
	end if;
	if (ll=37 and cc>=175 and cc<180) then grbp<="110";
	end if;
	if (cc=183 and ll=37) then grbp<="110";
	end if;
	if (ll=37 and cc>=183 and cc<185) then grbp<="110";
	end if;
	if (ll=37 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=191 and ll=37) then grbp<="110";
	end if;
	if (ll=37 and cc>=191 and cc<193) then grbp<="110";
	end if;
	if (cc=218 and ll=37) then grbp<="110";
	end if;
	if (cc=0 and ll=38) then grbp<="110";
	end if;
	if (ll=38 and cc>=0 and cc<12) then grbp<="110";
	end if;
	if (ll=38 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (ll=38 and cc>=175 and cc<180) then grbp<="110";
	end if;
	if (cc=186 and ll=38) then grbp<="110";
	end if;
	if (ll=38 and cc>=186 and cc<190) then grbp<="110";
	end if;
	if (cc=209 and ll=38) then grbp<="110";
	end if;
	if (cc=218 and ll=38) then grbp<="110";
	end if;
	if (cc=0 and ll=39) then grbp<="110";
	end if;
	if (ll=39 and cc>=0 and cc<8) then grbp<="110";
	end if;
	if (ll=39 and cc>=9 and cc<11) then grbp<="110";
	end if;
	if (ll=39 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=39 and cc>=175 and cc<180) then grbp<="110";
	end if;
	if (cc=186 and ll=39) then grbp<="110";
	end if;
	if (cc=189 and ll=39) then grbp<="110";
	end if;
	if (cc=209 and ll=39) then grbp<="110";
	end if;
	if (cc=219 and ll=39) then grbp<="110";
	end if;
	if (cc=0 and ll=40) then grbp<="110";
	end if;
	if (ll=40 and cc>=0 and cc<11) then grbp<="110";
	end if;
	if (ll=40 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=178 and ll=40) then grbp<="110";
	end if;
	if (cc=180 and ll=40) then grbp<="110";
	end if;
	if (cc=187 and ll=40) then grbp<="110";
	end if;
	if (cc=189 and ll=40) then grbp<="110";
	end if;
	if (cc=210 and ll=40) then grbp<="110";
	end if;
	if (cc=219 and ll=40) then grbp<="110";
	end if;
	if (cc=0 and ll=41) then grbp<="110";
	end if;
	if (ll=41 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (ll=41 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=186 and ll=41) then grbp<="110";
	end if;
	if (cc=188 and ll=41) then grbp<="110";
	end if;
	if (ll=41 and cc>=188 and cc<190) then grbp<="110";
	end if;
	if (cc=0 and ll=42) then grbp<="110";
	end if;
	if (ll=42 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (ll=42 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=179 and ll=42) then grbp<="110";
	end if;
	if (cc=181 and ll=42) then grbp<="110";
	end if;
	if (ll=42 and cc>=181 and cc<183) then grbp<="110";
	end if;
	if (cc=210 and ll=42) then grbp<="110";
	end if;
	if (cc=220 and ll=42) then grbp<="110";
	end if;
	if (cc=0 and ll=43) then grbp<="110";
	end if;
	if (ll=43 and cc>=0 and cc<9) then grbp<="110";
	end if;
	if (ll=43 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=43 and cc>=178 and cc<180) then grbp<="110";
	end if;
	if (cc=211 and ll=43) then grbp<="110";
	end if;
	if (cc=220 and ll=43) then grbp<="110";
	end if;
	if (cc=0 and ll=44) then grbp<="110";
	end if;
	if (ll=44 and cc>=0 and cc<9) then grbp<="110";
	end if;
	if (ll=44 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=0 and ll=45) then grbp<="110";
	end if;
	if (ll=45 and cc>=0 and cc<10) then grbp<="110";
	end if;
	if (ll=45 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=179 and ll=45) then grbp<="110";
	end if;
	if (cc=212 and ll=45) then grbp<="110";
	end if;
	if (cc=221 and ll=45) then grbp<="110";
	end if;
	if (cc=0 and ll=46) then grbp<="110";
	end if;
	if (ll=46 and cc>=0 and cc<9) then grbp<="110";
	end if;
	if (ll=46 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=0 and ll=47) then grbp<="110";
	end if;
	if (ll=47 and cc>=0 and cc<8) then grbp<="110";
	end if;
	if (ll=47 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=181 and ll=47) then grbp<="110";
	end if;
	if (cc=212 and ll=47) then grbp<="110";
	end if;
	if (cc=0 and ll=48) then grbp<="110";
	end if;
	if (ll=48 and cc>=0 and cc<8) then grbp<="110";
	end if;
	if (ll=48 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=181 and ll=48) then grbp<="110";
	end if;
	if (cc=222 and ll=48) then grbp<="110";
	end if;
	if (cc=0 and ll=49) then grbp<="110";
	end if;
	if (ll=49 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=49 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=213 and ll=49) then grbp<="110";
	end if;
	if (cc=222 and ll=49) then grbp<="110";
	end if;
	if (cc=0 and ll=50) then grbp<="110";
	end if;
	if (ll=50 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=50 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=83 and ll=50) then grbp<="110";
	end if;
	if (cc=104 and ll=50) then grbp<="110";
	end if;
	if (cc=213 and ll=50) then grbp<="110";
	end if;
	if (cc=222 and ll=50) then grbp<="110";
	end if;
	if (cc=0 and ll=51) then grbp<="110";
	end if;
	if (ll=51 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=51 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=52 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=52 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=109 and ll=52) then grbp<="110";
	end if;
	if (cc=183 and ll=52) then grbp<="110";
	end if;
	if (cc=214 and ll=52) then grbp<="110";
	end if;
	if (cc=221 and ll=52) then grbp<="110";
	end if;
	if (cc=0 and ll=53) then grbp<="110";
	end if;
	if (ll=53 and cc>=0 and cc<7) then grbp<="110";
	end if;
	if (ll=53 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (ll=53 and cc>=77 and cc<79) then grbp<="110";
	end if;
	if (cc=214 and ll=53) then grbp<="110";
	end if;
	if (cc=221 and ll=53) then grbp<="110";
	end if;
	if (cc=0 and ll=54) then grbp<="110";
	end if;
	if (ll=54 and cc>=0 and cc<6) then grbp<="110";
	end if;
	if (ll=54 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=215 and ll=54) then grbp<="110";
	end if;
	if (cc=220 and ll=54) then grbp<="110";
	end if;
	if (cc=0 and ll=55) then grbp<="110";
	end if;
	if (ll=55 and cc>=0 and cc<6) then grbp<="110";
	end if;
	if (ll=55 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=220 and ll=55) then grbp<="110";
	end if;
	if (cc=0 and ll=56) then grbp<="110";
	end if;
	if (ll=56 and cc>=0 and cc<5) then grbp<="110";
	end if;
	if (ll=56 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=215 and ll=56) then grbp<="110";
	end if;
	if (cc=219 and ll=56) then grbp<="110";
	end if;
	if (cc=0 and ll=57) then grbp<="110";
	end if;
	if (ll=57 and cc>=0 and cc<5) then grbp<="110";
	end if;
	if (ll=57 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=109 and ll=57) then grbp<="110";
	end if;
	if (cc=0 and ll=58) then grbp<="110";
	end if;
	if (ll=58 and cc>=0 and cc<5) then grbp<="110";
	end if;
	if (ll=58 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=218 and ll=58) then grbp<="110";
	end if;
	if (cc=0 and ll=59) then grbp<="110";
	end if;
	if (ll=59 and cc>=0 and cc<5) then grbp<="110";
	end if;
	if (ll=59 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=216 and ll=59) then grbp<="110";
	end if;
	if (ll=59 and cc>=216 and cc<218) then grbp<="110";
	end if;
	if (ll=60 and cc>=0 and cc<4) then grbp<="110";
	end if;
	if (ll=60 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (ll=60 and cc>=214 and cc<217) then grbp<="110";
	end if;
	if (ll=61 and cc>=0 and cc<4) then grbp<="110";
	end if;
	if (ll=61 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=0 and ll=62) then grbp<="110";
	end if;
	if (ll=62 and cc>=0 and cc<4) then grbp<="110";
	end if;
	if (ll=62 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=108 and ll=62) then grbp<="110";
	end if;
	if (ll=62 and cc>=108 and cc<110) then grbp<="110";
	end if;
	if (ll=62 and cc>=170 and cc<172) then grbp<="110";
	end if;
	if (ll=63 and cc>=1 and cc<3) then grbp<="110";
	end if;
	if (ll=63 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=106 and ll=63) then grbp<="110";
	end if;
	if (cc=108 and ll=63) then grbp<="110";
	end if;
	if (cc=111 and ll=63) then grbp<="110";
	end if;
	if (cc=168 and ll=63) then grbp<="110";
	end if;
	if (ll=63 and cc>=168 and cc<170) then grbp<="110";
	end if;
	if (ll=63 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=0 and ll=64) then grbp<="110";
	end if;
	if (ll=64 and cc>=0 and cc<3) then grbp<="110";
	end if;
	if (ll=64 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=168 and ll=64) then grbp<="110";
	end if;
	if (cc=170 and ll=64) then grbp<="110";
	end if;
	if (cc=213 and ll=64) then grbp<="110";
	end if;
	if (ll=64 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=0 and ll=65) then grbp<="110";
	end if;
	if (ll=65 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=65 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=212 and ll=65) then grbp<="110";
	end if;
	if (ll=65 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=0 and ll=66) then grbp<="110";
	end if;
	if (ll=66 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=66 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=169 and ll=66) then grbp<="110";
	end if;
	if (cc=212 and ll=66) then grbp<="110";
	end if;
	if (cc=249 and ll=66) then grbp<="110";
	end if;
	if (ll=66 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=67 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=67 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (ll=67 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=68 and cc>=0 and cc<2) then grbp<="110";
	end if;
	if (ll=68 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=211 and ll=68) then grbp<="110";
	end if;
	if (ll=68 and cc>=211 and cc<213) then grbp<="110";
	end if;
	if (ll=68 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (cc=17 and ll=69) then grbp<="110";
	end if;
	if (ll=69 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=110 and ll=69) then grbp<="110";
	end if;
	if (cc=169 and ll=69) then grbp<="110";
	end if;
	if (cc=249 and ll=69) then grbp<="110";
	end if;
	if (ll=69 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=70 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=250 and ll=70) then grbp<="110";
	end if;
	if (cc=17 and ll=71) then grbp<="110";
	end if;
	if (ll=71 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=247 and ll=71) then grbp<="110";
	end if;
	if (cc=250 and ll=71) then grbp<="110";
	end if;
	if (cc=17 and ll=72) then grbp<="110";
	end if;
	if (ll=72 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=16 and ll=73) then grbp<="110";
	end if;
	if (ll=73 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (ll=73 and cc>=107 and cc<111) then grbp<="110";
	end if;
	if (cc=247 and ll=73) then grbp<="110";
	end if;
	if (cc=17 and ll=74) then grbp<="110";
	end if;
	if (ll=74 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=246 and ll=74) then grbp<="110";
	end if;
	if (ll=74 and cc>=246 and cc<248) then grbp<="110";
	end if;
	if (ll=75 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=170 and ll=75) then grbp<="110";
	end if;
	if (cc=246 and ll=75) then grbp<="110";
	end if;
	if (ll=75 and cc>=246 and cc<248) then grbp<="110";
	end if;
	if (cc=17 and ll=76) then grbp<="110";
	end if;
	if (ll=76 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=246 and ll=76) then grbp<="110";
	end if;
	if (ll=76 and cc>=246 and cc<248) then grbp<="110";
	end if;
	if (cc=16 and ll=77) then grbp<="110";
	end if;
	if (ll=77 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=246 and ll=77) then grbp<="110";
	end if;
	if (cc=249 and ll=77) then grbp<="110";
	end if;
	if (ll=77 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=78 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=78 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=79 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=116 and ll=79) then grbp<="110";
	end if;
	if (cc=248 and ll=79) then grbp<="110";
	end if;
	if (ll=79 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=80 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=114 and ll=80) then grbp<="110";
	end if;
	if (cc=248 and ll=80) then grbp<="110";
	end if;
	if (ll=80 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=81 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=113 and ll=81) then grbp<="110";
	end if;
	if (cc=168 and ll=81) then grbp<="110";
	end if;
	if (cc=171 and ll=81) then grbp<="110";
	end if;
	if (cc=244 and ll=81) then grbp<="110";
	end if;
	if (cc=247 and ll=81) then grbp<="110";
	end if;
	if (ll=81 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=82 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=175 and ll=82) then grbp<="110";
	end if;
	if (cc=244 and ll=82) then grbp<="110";
	end if;
	if (cc=247 and ll=82) then grbp<="110";
	end if;
	if (cc=17 and ll=83) then grbp<="110";
	end if;
	if (ll=83 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=168 and ll=83) then grbp<="110";
	end if;
	if (cc=243 and ll=83) then grbp<="110";
	end if;
	if (cc=246 and ll=83) then grbp<="110";
	end if;
	if (ll=83 and cc>=246 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=84) then grbp<="110";
	end if;
	if (ll=84 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=249 and ll=84) then grbp<="110";
	end if;
	if (ll=84 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=85 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=245 and ll=85) then grbp<="110";
	end if;
	if (ll=85 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (cc=17 and ll=86) then grbp<="110";
	end if;
	if (ll=86 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=86 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (cc=17 and ll=87) then grbp<="110";
	end if;
	if (ll=87 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=249 and ll=87) then grbp<="110";
	end if;
	if (cc=17 and ll=88) then grbp<="110";
	end if;
	if (ll=88 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=244 and ll=88) then grbp<="110";
	end if;
	if (cc=247 and ll=88) then grbp<="110";
	end if;
	if (cc=249 and ll=88) then grbp<="110";
	end if;
	if (ll=88 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=89 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=243 and ll=89) then grbp<="110";
	end if;
	if (ll=89 and cc>=243 and cc<248) then grbp<="110";
	end if;
	if (ll=89 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=90 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=244 and ll=90) then grbp<="110";
	end if;
	if (cc=246 and ll=90) then grbp<="110";
	end if;
	if (ll=90 and cc>=246 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=91) then grbp<="110";
	end if;
	if (ll=91 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=242 and ll=91) then grbp<="110";
	end if;
	if (ll=91 and cc>=242 and cc<251) then grbp<="110";
	end if;
	if (ll=92 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=92 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=245 and ll=92) then grbp<="110";
	end if;
	if (cc=249 and ll=92) then grbp<="110";
	end if;
	if (ll=92 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=93 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=174 and ll=93) then grbp<="110";
	end if;
	if (ll=93 and cc>=174 and cc<176) then grbp<="110";
	end if;
	if (cc=243 and ll=93) then grbp<="110";
	end if;
	if (cc=246 and ll=93) then grbp<="110";
	end if;
	if (ll=93 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=94 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=243 and ll=94) then grbp<="110";
	end if;
	if (ll=94 and cc>=243 and cc<245) then grbp<="110";
	end if;
	if (ll=94 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=95 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=106 and ll=95) then grbp<="110";
	end if;
	if (cc=235 and ll=95) then grbp<="110";
	end if;
	if (cc=243 and ll=95) then grbp<="110";
	end if;
	if (ll=95 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=96 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=240 and ll=96) then grbp<="110";
	end if;
	if (cc=243 and ll=96) then grbp<="110";
	end if;
	if (ll=96 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=97 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=239 and ll=97) then grbp<="110";
	end if;
	if (ll=97 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=97 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=98 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=239 and ll=98) then grbp<="110";
	end if;
	if (cc=243 and ll=98) then grbp<="110";
	end if;
	if (cc=245 and ll=98) then grbp<="110";
	end if;
	if (ll=98 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=99 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=234 and ll=99) then grbp<="110";
	end if;
	if (cc=239 and ll=99) then grbp<="110";
	end if;
	if (cc=243 and ll=99) then grbp<="110";
	end if;
	if (ll=99 and cc>=243 and cc<245) then grbp<="110";
	end if;
	if (ll=99 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=100 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=100 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=233 and ll=100) then grbp<="110";
	end if;
	if (cc=239 and ll=100) then grbp<="110";
	end if;
	if (cc=242 and ll=100) then grbp<="110";
	end if;
	if (cc=244 and ll=100) then grbp<="110";
	end if;
	if (cc=247 and ll=100) then grbp<="110";
	end if;
	if (ll=100 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=101 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=63 and ll=101) then grbp<="110";
	end if;
	if (cc=107 and ll=101) then grbp<="110";
	end if;
	if (cc=168 and ll=101) then grbp<="110";
	end if;
	if (cc=170 and ll=101) then grbp<="110";
	end if;
	if (cc=233 and ll=101) then grbp<="110";
	end if;
	if (cc=239 and ll=101) then grbp<="110";
	end if;
	if (ll=101 and cc>=239 and cc<243) then grbp<="110";
	end if;
	if (ll=101 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (ll=101 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=102 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=168 and ll=102) then grbp<="110";
	end if;
	if (cc=171 and ll=102) then grbp<="110";
	end if;
	if (cc=232 and ll=102) then grbp<="110";
	end if;
	if (cc=243 and ll=102) then grbp<="110";
	end if;
	if (ll=102 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=103 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=168 and ll=103) then grbp<="110";
	end if;
	if (ll=103 and cc>=168 and cc<170) then grbp<="110";
	end if;
	if (ll=103 and cc>=171 and cc<175) then grbp<="110";
	end if;
	if (cc=240 and ll=103) then grbp<="110";
	end if;
	if (ll=103 and cc>=240 and cc<246) then grbp<="110";
	end if;
	if (ll=103 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=104 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=104 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (ll=104 and cc>=171 and cc<173) then grbp<="110";
	end if;
	if (cc=189 and ll=104) then grbp<="110";
	end if;
	if (cc=238 and ll=104) then grbp<="110";
	end if;
	if (ll=104 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=105 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=171 and ll=105) then grbp<="110";
	end if;
	if (cc=174 and ll=105) then grbp<="110";
	end if;
	if (cc=238 and ll=105) then grbp<="110";
	end if;
	if (ll=105 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=106 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=106 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (cc=171 and ll=106) then grbp<="110";
	end if;
	if (cc=173 and ll=106) then grbp<="110";
	end if;
	if (cc=235 and ll=106) then grbp<="110";
	end if;
	if (cc=237 and ll=106) then grbp<="110";
	end if;
	if (cc=239 and ll=106) then grbp<="110";
	end if;
	if (ll=106 and cc>=239 and cc<243) then grbp<="110";
	end if;
	if (cc=246 and ll=106) then grbp<="110";
	end if;
	if (ll=106 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=107 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=107 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (cc=231 and ll=107) then grbp<="110";
	end if;
	if (cc=236 and ll=107) then grbp<="110";
	end if;
	if (ll=107 and cc>=236 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=108) then grbp<="110";
	end if;
	if (ll=108 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=62 and ll=108) then grbp<="110";
	end if;
	if (ll=108 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (cc=105 and ll=108) then grbp<="110";
	end if;
	if (ll=108 and cc>=105 and cc<107) then grbp<="110";
	end if;
	if (cc=234 and ll=108) then grbp<="110";
	end if;
	if (cc=236 and ll=108) then grbp<="110";
	end if;
	if (cc=239 and ll=108) then grbp<="110";
	end if;
	if (ll=108 and cc>=239 and cc<246) then grbp<="110";
	end if;
	if (ll=108 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=109 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=172 and ll=109) then grbp<="110";
	end if;
	if (cc=230 and ll=109) then grbp<="110";
	end if;
	if (cc=234 and ll=109) then grbp<="110";
	end if;
	if (ll=109 and cc>=234 and cc<237) then grbp<="110";
	end if;
	if (cc=240 and ll=109) then grbp<="110";
	end if;
	if (ll=109 and cc>=240 and cc<251) then grbp<="110";
	end if;
	if (ll=110 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=94 and ll=110) then grbp<="110";
	end if;
	if (cc=96 and ll=110) then grbp<="110";
	end if;
	if (ll=110 and cc>=96 and cc<98) then grbp<="110";
	end if;
	if (cc=238 and ll=110) then grbp<="110";
	end if;
	if (ll=110 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=111 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=94 and ll=111) then grbp<="110";
	end if;
	if (cc=98 and ll=111) then grbp<="110";
	end if;
	if (cc=233 and ll=111) then grbp<="110";
	end if;
	if (cc=238 and ll=111) then grbp<="110";
	end if;
	if (ll=111 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=111 and cc>=241 and cc<250) then grbp<="110";
	end if;
	if (ll=112 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=93 and ll=112) then grbp<="110";
	end if;
	if (ll=112 and cc>=93 and cc<97) then grbp<="110";
	end if;
	if (cc=169 and ll=112) then grbp<="110";
	end if;
	if (cc=228 and ll=112) then grbp<="110";
	end if;
	if (cc=233 and ll=112) then grbp<="110";
	end if;
	if (ll=112 and cc>=233 and cc<243) then grbp<="110";
	end if;
	if (cc=246 and ll=112) then grbp<="110";
	end if;
	if (ll=112 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=113 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=95 and ll=113) then grbp<="110";
	end if;
	if (cc=234 and ll=113) then grbp<="110";
	end if;
	if (ll=113 and cc>=234 and cc<238) then grbp<="110";
	end if;
	if (ll=113 and cc>=240 and cc<251) then grbp<="110";
	end if;
	if (ll=114 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=92 and ll=114) then grbp<="110";
	end if;
	if (ll=114 and cc>=92 and cc<94) then grbp<="110";
	end if;
	if (cc=232 and ll=114) then grbp<="110";
	end if;
	if (ll=114 and cc>=232 and cc<240) then grbp<="110";
	end if;
	if (ll=114 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=115 and cc>=18 and cc<27) then grbp<="110";
	end if;
	if (cc=93 and ll=115) then grbp<="110";
	end if;
	if (cc=99 and ll=115) then grbp<="110";
	end if;
	if (cc=227 and ll=115) then grbp<="110";
	end if;
	if (ll=115 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=115 and cc>=232 and cc<237) then grbp<="110";
	end if;
	if (ll=115 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=116 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=116 and cc>=93 and cc<95) then grbp<="110";
	end if;
	if (cc=232 and ll=116) then grbp<="110";
	end if;
	if (ll=116 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (cc=238 and ll=116) then grbp<="110";
	end if;
	if (ll=116 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=117 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=117) then grbp<="110";
	end if;
	if (ll=117 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=93 and ll=117) then grbp<="110";
	end if;
	if (cc=227 and ll=117) then grbp<="110";
	end if;
	if (cc=231 and ll=117) then grbp<="110";
	end if;
	if (ll=117 and cc>=231 and cc<234) then grbp<="110";
	end if;
	if (ll=117 and cc>=235 and cc<246) then grbp<="110";
	end if;
	if (ll=117 and cc>=247 and cc<250) then grbp<="110";
	end if;
	if (ll=118 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=118 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=238 and ll=118) then grbp<="110";
	end if;
	if (ll=118 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (cc=243 and ll=118) then grbp<="110";
	end if;
	if (ll=118 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=119 and cc>=16 and cc<24) then grbp<="110";
	end if;
	if (ll=119 and cc>=25 and cc<28) then grbp<="110";
	end if;
	if (cc=96 and ll=119) then grbp<="110";
	end if;
	if (cc=99 and ll=119) then grbp<="110";
	end if;
	if (cc=106 and ll=119) then grbp<="110";
	end if;
	if (cc=232 and ll=119) then grbp<="110";
	end if;
	if (ll=119 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (ll=119 and cc>=237 and cc<240) then grbp<="110";
	end if;
	if (ll=119 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=120 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=120 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=115 and ll=120) then grbp<="110";
	end if;
	if (ll=120 and cc>=115 and cc<117) then grbp<="110";
	end if;
	if (cc=233 and ll=120) then grbp<="110";
	end if;
	if (ll=120 and cc>=233 and cc<236) then grbp<="110";
	end if;
	if (ll=120 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=121 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=121 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=233 and ll=121) then grbp<="110";
	end if;
	if (ll=121 and cc>=233 and cc<237) then grbp<="110";
	end if;
	if (ll=121 and cc>=239 and cc<251) then grbp<="110";
	end if;
	if (ll=122 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=122 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=99 and ll=122) then grbp<="110";
	end if;
	if (cc=103 and ll=122) then grbp<="110";
	end if;
	if (ll=122 and cc>=103 and cc<106) then grbp<="110";
	end if;
	if (cc=225 and ll=122) then grbp<="110";
	end if;
	if (cc=231 and ll=122) then grbp<="110";
	end if;
	if (ll=122 and cc>=231 and cc<234) then grbp<="110";
	end if;
	if (cc=237 and ll=122) then grbp<="110";
	end if;
	if (cc=239 and ll=122) then grbp<="110";
	end if;
	if (ll=122 and cc>=239 and cc<251) then grbp<="110";
	end if;
	if (ll=123 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=93 and ll=123) then grbp<="110";
	end if;
	if (cc=99 and ll=123) then grbp<="110";
	end if;
	if (cc=101 and ll=123) then grbp<="110";
	end if;
	if (cc=237 and ll=123) then grbp<="110";
	end if;
	if (cc=239 and ll=123) then grbp<="110";
	end if;
	if (ll=123 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=123 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (ll=123 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=124 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=124 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=92 and ll=124) then grbp<="110";
	end if;
	if (cc=102 and ll=124) then grbp<="110";
	end if;
	if (cc=229 and ll=124) then grbp<="110";
	end if;
	if (cc=232 and ll=124) then grbp<="110";
	end if;
	if (ll=124 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (ll=124 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (ll=124 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (cc=245 and ll=124) then grbp<="110";
	end if;
	if (ll=124 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=125 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=125 and cc>=60 and cc<64) then grbp<="110";
	end if;
	if (cc=111 and ll=125) then grbp<="110";
	end if;
	if (ll=125 and cc>=111 and cc<113) then grbp<="110";
	end if;
	if (cc=232 and ll=125) then grbp<="110";
	end if;
	if (ll=125 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (cc=237 and ll=125) then grbp<="110";
	end if;
	if (cc=239 and ll=125) then grbp<="110";
	end if;
	if (ll=125 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (cc=245 and ll=125) then grbp<="110";
	end if;
	if (ll=125 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=126 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=126 and cc>=60 and cc<62) then grbp<="110";
	end if;
	if (cc=117 and ll=126) then grbp<="110";
	end if;
	if (cc=230 and ll=126) then grbp<="110";
	end if;
	if (ll=126 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=126 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (ll=126 and cc>=239 and cc<251) then grbp<="110";
	end if;
	if (ll=127 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=127 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (ll=127 and cc>=98 and cc<100) then grbp<="110";
	end if;
	if (cc=106 and ll=127) then grbp<="110";
	end if;
	if (cc=118 and ll=127) then grbp<="110";
	end if;
	if (cc=130 and ll=127) then grbp<="110";
	end if;
	if (cc=223 and ll=127) then grbp<="110";
	end if;
	if (cc=230 and ll=127) then grbp<="110";
	end if;
	if (ll=127 and cc>=230 and cc<233) then grbp<="110";
	end if;
	if (ll=127 and cc>=234 and cc<236) then grbp<="110";
	end if;
	if (cc=239 and ll=127) then grbp<="110";
	end if;
	if (cc=241 and ll=127) then grbp<="110";
	end if;
	if (ll=127 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=128 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=128 and cc>=60 and cc<63) then grbp<="110";
	end if;
	if (cc=97 and ll=128) then grbp<="110";
	end if;
	if (ll=128 and cc>=97 and cc<99) then grbp<="110";
	end if;
	if (cc=230 and ll=128) then grbp<="110";
	end if;
	if (cc=233 and ll=128) then grbp<="110";
	end if;
	if (ll=128 and cc>=233 and cc<235) then grbp<="110";
	end if;
	if (ll=128 and cc>=237 and cc<251) then grbp<="110";
	end if;
	if (ll=129 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (ll=129 and cc>=60 and cc<65) then grbp<="110";
	end if;
	if (cc=238 and ll=129) then grbp<="110";
	end if;
	if (ll=129 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=130 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=130 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (cc=89 and ll=130) then grbp<="110";
	end if;
	if (cc=103 and ll=130) then grbp<="110";
	end if;
	if (cc=124 and ll=130) then grbp<="110";
	end if;
	if (cc=132 and ll=130) then grbp<="110";
	end if;
	if (cc=231 and ll=130) then grbp<="110";
	end if;
	if (cc=233 and ll=130) then grbp<="110";
	end if;
	if (cc=235 and ll=130) then grbp<="110";
	end if;
	if (cc=237 and ll=130) then grbp<="110";
	end if;
	if (ll=130 and cc>=237 and cc<249) then grbp<="110";
	end if;
	if (cc=16 and ll=131) then grbp<="110";
	end if;
	if (ll=131 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=62 and ll=131) then grbp<="110";
	end if;
	if (ll=131 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (ll=131 and cc>=106 and cc<108) then grbp<="110";
	end if;
	if (cc=229 and ll=131) then grbp<="110";
	end if;
	if (cc=231 and ll=131) then grbp<="110";
	end if;
	if (ll=131 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (cc=239 and ll=131) then grbp<="110";
	end if;
	if (cc=241 and ll=131) then grbp<="110";
	end if;
	if (cc=243 and ll=131) then grbp<="110";
	end if;
	if (ll=131 and cc>=243 and cc<245) then grbp<="110";
	end if;
	if (cc=248 and ll=131) then grbp<="110";
	end if;
	if (ll=131 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=132 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=132 and cc>=60 and cc<62) then grbp<="110";
	end if;
	if (ll=132 and cc>=63 and cc<66) then grbp<="110";
	end if;
	if (cc=100 and ll=132) then grbp<="110";
	end if;
	if (cc=104 and ll=132) then grbp<="110";
	end if;
	if (cc=109 and ll=132) then grbp<="110";
	end if;
	if (cc=122 and ll=132) then grbp<="110";
	end if;
	if (cc=155 and ll=132) then grbp<="110";
	end if;
	if (cc=237 and ll=132) then grbp<="110";
	end if;
	if (ll=132 and cc>=237 and cc<241) then grbp<="110";
	end if;
	if (ll=132 and cc>=242 and cc<250) then grbp<="110";
	end if;
	if (ll=133 and cc>=17 and cc<27) then grbp<="110";
	end if;
	if (cc=61 and ll=133) then grbp<="110";
	end if;
	if (ll=133 and cc>=61 and cc<66) then grbp<="110";
	end if;
	if (cc=99 and ll=133) then grbp<="110";
	end if;
	if (cc=228 and ll=133) then grbp<="110";
	end if;
	if (cc=232 and ll=133) then grbp<="110";
	end if;
	if (cc=234 and ll=133) then grbp<="110";
	end if;
	if (ll=133 and cc>=234 and cc<251) then grbp<="110";
	end if;
	if (ll=134 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=60 and ll=134) then grbp<="110";
	end if;
	if (ll=134 and cc>=60 and cc<65) then grbp<="110";
	end if;
	if (cc=107 and ll=134) then grbp<="110";
	end if;
	if (cc=123 and ll=134) then grbp<="110";
	end if;
	if (cc=127 and ll=134) then grbp<="110";
	end if;
	if (ll=134 and cc>=127 and cc<129) then grbp<="110";
	end if;
	if (cc=194 and ll=134) then grbp<="110";
	end if;
	if (cc=221 and ll=134) then grbp<="110";
	end if;
	if (cc=232 and ll=134) then grbp<="110";
	end if;
	if (ll=134 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (cc=238 and ll=134) then grbp<="110";
	end if;
	if (ll=134 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=135 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=135 and cc>=60 and cc<64) then grbp<="110";
	end if;
	if (cc=108 and ll=135) then grbp<="110";
	end if;
	if (cc=112 and ll=135) then grbp<="110";
	end if;
	if (cc=114 and ll=135) then grbp<="110";
	end if;
	if (cc=117 and ll=135) then grbp<="110";
	end if;
	if (ll=135 and cc>=117 and cc<119) then grbp<="110";
	end if;
	if (cc=225 and ll=135) then grbp<="110";
	end if;
	if (cc=227 and ll=135) then grbp<="110";
	end if;
	if (cc=232 and ll=135) then grbp<="110";
	end if;
	if (ll=135 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (ll=135 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (ll=135 and cc>=239 and cc<247) then grbp<="110";
	end if;
	if (ll=135 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=136 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=136 and cc>=59 and cc<64) then grbp<="110";
	end if;
	if (cc=102 and ll=136) then grbp<="110";
	end if;
	if (cc=124 and ll=136) then grbp<="110";
	end if;
	if (ll=136 and cc>=124 and cc<126) then grbp<="110";
	end if;
	if (cc=193 and ll=136) then grbp<="110";
	end if;
	if (cc=227 and ll=136) then grbp<="110";
	end if;
	if (ll=136 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=136 and cc>=230 and cc<235) then grbp<="110";
	end if;
	if (ll=136 and cc>=237 and cc<239) then grbp<="110";
	end if;
	if (ll=136 and cc>=240 and cc<251) then grbp<="110";
	end if;
	if (ll=137 and cc>=16 and cc<27) then grbp<="110";
	end if;
	if (cc=61 and ll=137) then grbp<="110";
	end if;
	if (ll=137 and cc>=61 and cc<64) then grbp<="110";
	end if;
	if (cc=92 and ll=137) then grbp<="110";
	end if;
	if (cc=100 and ll=137) then grbp<="110";
	end if;
	if (cc=105 and ll=137) then grbp<="110";
	end if;
	if (cc=227 and ll=137) then grbp<="110";
	end if;
	if (ll=137 and cc>=227 and cc<230) then grbp<="110";
	end if;
	if (ll=137 and cc>=233 and cc<236) then grbp<="110";
	end if;
	if (cc=239 and ll=137) then grbp<="110";
	end if;
	if (cc=241 and ll=137) then grbp<="110";
	end if;
	if (ll=137 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=138 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=138 and cc>=60 and cc<65) then grbp<="110";
	end if;
	if (cc=105 and ll=138) then grbp<="110";
	end if;
	if (cc=107 and ll=138) then grbp<="110";
	end if;
	if (cc=230 and ll=138) then grbp<="110";
	end if;
	if (cc=232 and ll=138) then grbp<="110";
	end if;
	if (ll=138 and cc>=232 and cc<236) then grbp<="110";
	end if;
	if (cc=239 and ll=138) then grbp<="110";
	end if;
	if (ll=138 and cc>=239 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=139) then grbp<="110";
	end if;
	if (ll=139 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=139 and cc>=60 and cc<66) then grbp<="110";
	end if;
	if (cc=106 and ll=139) then grbp<="110";
	end if;
	if (ll=139 and cc>=106 and cc<108) then grbp<="110";
	end if;
	if (cc=138 and ll=139) then grbp<="110";
	end if;
	if (cc=191 and ll=139) then grbp<="110";
	end if;
	if (cc=224 and ll=139) then grbp<="110";
	end if;
	if (ll=139 and cc>=224 and cc<236) then grbp<="110";
	end if;
	if (ll=139 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=139 and cc>=242 and cc<251) then grbp<="110";
	end if;
	if (ll=140 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=63 and ll=140) then grbp<="110";
	end if;
	if (cc=65 and ll=140) then grbp<="110";
	end if;
	if (ll=140 and cc>=65 and cc<67) then grbp<="110";
	end if;
	if (cc=124 and ll=140) then grbp<="110";
	end if;
	if (cc=130 and ll=140) then grbp<="110";
	end if;
	if (cc=193 and ll=140) then grbp<="110";
	end if;
	if (cc=223 and ll=140) then grbp<="110";
	end if;
	if (cc=225 and ll=140) then grbp<="110";
	end if;
	if (ll=140 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=140 and cc>=228 and cc<237) then grbp<="110";
	end if;
	if (ll=140 and cc>=238 and cc<247) then grbp<="110";
	end if;
	if (ll=140 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=141 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=141 and cc>=60 and cc<62) then grbp<="110";
	end if;
	if (ll=141 and cc>=64 and cc<67) then grbp<="110";
	end if;
	if (cc=104 and ll=141) then grbp<="110";
	end if;
	if (cc=125 and ll=141) then grbp<="110";
	end if;
	if (cc=128 and ll=141) then grbp<="110";
	end if;
	if (ll=141 and cc>=128 and cc<130) then grbp<="110";
	end if;
	if (cc=218 and ll=141) then grbp<="110";
	end if;
	if (cc=224 and ll=141) then grbp<="110";
	end if;
	if (cc=226 and ll=141) then grbp<="110";
	end if;
	if (ll=141 and cc>=226 and cc<232) then grbp<="110";
	end if;
	if (ll=141 and cc>=233 and cc<248) then grbp<="110";
	end if;
	if (ll=141 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=142 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=142 and cc>=60 and cc<63) then grbp<="110";
	end if;
	if (cc=66 and ll=142) then grbp<="110";
	end if;
	if (cc=105 and ll=142) then grbp<="110";
	end if;
	if (cc=144 and ll=142) then grbp<="110";
	end if;
	if (cc=187 and ll=142) then grbp<="110";
	end if;
	if (cc=189 and ll=142) then grbp<="110";
	end if;
	if (cc=218 and ll=142) then grbp<="110";
	end if;
	if (cc=223 and ll=142) then grbp<="110";
	end if;
	if (cc=225 and ll=142) then grbp<="110";
	end if;
	if (ll=142 and cc>=225 and cc<229) then grbp<="110";
	end if;
	if (ll=142 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (cc=239 and ll=142) then grbp<="110";
	end if;
	if (ll=142 and cc>=239 and cc<251) then grbp<="110";
	end if;
	if (ll=143 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=143 and cc>=61 and cc<64) then grbp<="110";
	end if;
	if (cc=67 and ll=143) then grbp<="110";
	end if;
	if (cc=189 and ll=143) then grbp<="110";
	end if;
	if (cc=222 and ll=143) then grbp<="110";
	end if;
	if (ll=143 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=143 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (ll=143 and cc>=229 and cc<235) then grbp<="110";
	end if;
	if (ll=143 and cc>=236 and cc<251) then grbp<="110";
	end if;
	if (ll=144 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=63 and ll=144) then grbp<="110";
	end if;
	if (ll=144 and cc>=63 and cc<68) then grbp<="110";
	end if;
	if (cc=222 and ll=144) then grbp<="110";
	end if;
	if (cc=225 and ll=144) then grbp<="110";
	end if;
	if (cc=227 and ll=144) then grbp<="110";
	end if;
	if (ll=144 and cc>=227 and cc<232) then grbp<="110";
	end if;
	if (ll=144 and cc>=233 and cc<240) then grbp<="110";
	end if;
	if (ll=144 and cc>=241 and cc<245) then grbp<="110";
	end if;
	if (ll=144 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=145 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=63 and ll=145) then grbp<="110";
	end if;
	if (ll=145 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=68 and ll=145) then grbp<="110";
	end if;
	if (cc=70 and ll=145) then grbp<="110";
	end if;
	if (cc=149 and ll=145) then grbp<="110";
	end if;
	if (cc=225 and ll=145) then grbp<="110";
	end if;
	if (cc=228 and ll=145) then grbp<="110";
	end if;
	if (ll=145 and cc>=228 and cc<233) then grbp<="110";
	end if;
	if (cc=238 and ll=145) then grbp<="110";
	end if;
	if (ll=145 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=146 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=62 and ll=146) then grbp<="110";
	end if;
	if (cc=64 and ll=146) then grbp<="110";
	end if;
	if (ll=146 and cc>=64 and cc<66) then grbp<="110";
	end if;
	if (cc=186 and ll=146) then grbp<="110";
	end if;
	if (cc=226 and ll=146) then grbp<="110";
	end if;
	if (ll=146 and cc>=226 and cc<250) then grbp<="110";
	end if;
	if (ll=147 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=147) then grbp<="110";
	end if;
	if (cc=63 and ll=147) then grbp<="110";
	end if;
	if (ll=147 and cc>=63 and cc<66) then grbp<="110";
	end if;
	if (cc=69 and ll=147) then grbp<="110";
	end if;
	if (cc=71 and ll=147) then grbp<="110";
	end if;
	if (cc=147 and ll=147) then grbp<="110";
	end if;
	if (cc=185 and ll=147) then grbp<="110";
	end if;
	if (cc=225 and ll=147) then grbp<="110";
	end if;
	if (cc=229 and ll=147) then grbp<="110";
	end if;
	if (ll=147 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (cc=234 and ll=147) then grbp<="110";
	end if;
	if (ll=147 and cc>=234 and cc<237) then grbp<="110";
	end if;
	if (cc=240 and ll=147) then grbp<="110";
	end if;
	if (ll=147 and cc>=240 and cc<251) then grbp<="110";
	end if;
	if (ll=148 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=63 and ll=148) then grbp<="110";
	end if;
	if (cc=65 and ll=148) then grbp<="110";
	end if;
	if (ll=148 and cc>=65 and cc<67) then grbp<="110";
	end if;
	if (cc=146 and ll=148) then grbp<="110";
	end if;
	if (ll=148 and cc>=146 and cc<148) then grbp<="110";
	end if;
	if (cc=217 and ll=148) then grbp<="110";
	end if;
	if (cc=228 and ll=148) then grbp<="110";
	end if;
	if (ll=148 and cc>=228 and cc<230) then grbp<="110";
	end if;
	if (ll=148 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (cc=237 and ll=148) then grbp<="110";
	end if;
	if (ll=148 and cc>=237 and cc<251) then grbp<="110";
	end if;
	if (ll=149 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=62 and ll=149) then grbp<="110";
	end if;
	if (cc=64 and ll=149) then grbp<="110";
	end if;
	if (ll=149 and cc>=64 and cc<67) then grbp<="110";
	end if;
	if (cc=182 and ll=149) then grbp<="110";
	end if;
	if (cc=224 and ll=149) then grbp<="110";
	end if;
	if (cc=227 and ll=149) then grbp<="110";
	end if;
	if (ll=149 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (cc=232 and ll=149) then grbp<="110";
	end if;
	if (cc=234 and ll=149) then grbp<="110";
	end if;
	if (cc=236 and ll=149) then grbp<="110";
	end if;
	if (ll=149 and cc>=236 and cc<251) then grbp<="110";
	end if;
	if (ll=150 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=150) then grbp<="110";
	end if;
	if (ll=150 and cc>=61 and cc<63) then grbp<="110";
	end if;
	if (ll=150 and cc>=64 and cc<66) then grbp<="110";
	end if;
	if (ll=150 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (cc=236 and ll=150) then grbp<="110";
	end if;
	if (ll=150 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (ll=150 and cc>=239 and cc<251) then grbp<="110";
	end if;
	if (ll=151 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=151) then grbp<="110";
	end if;
	if (cc=63 and ll=151) then grbp<="110";
	end if;
	if (cc=65 and ll=151) then grbp<="110";
	end if;
	if (cc=179 and ll=151) then grbp<="110";
	end if;
	if (cc=196 and ll=151) then grbp<="110";
	end if;
	if (cc=224 and ll=151) then grbp<="110";
	end if;
	if (ll=151 and cc>=224 and cc<227) then grbp<="110";
	end if;
	if (cc=236 and ll=151) then grbp<="110";
	end if;
	if (ll=151 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (ll=151 and cc>=239 and cc<245) then grbp<="110";
	end if;
	if (ll=151 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=152 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=65 and ll=152) then grbp<="110";
	end if;
	if (ll=152 and cc>=65 and cc<67) then grbp<="110";
	end if;
	if (cc=178 and ll=152) then grbp<="110";
	end if;
	if (cc=195 and ll=152) then grbp<="110";
	end if;
	if (cc=223 and ll=152) then grbp<="110";
	end if;
	if (cc=225 and ll=152) then grbp<="110";
	end if;
	if (ll=152 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=152 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=152 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=152 and cc>=242 and cc<244) then grbp<="110";
	end if;
	if (ll=152 and cc>=245 and cc<248) then grbp<="110";
	end if;
	if (ll=152 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=153 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=64 and ll=153) then grbp<="110";
	end if;
	if (ll=153 and cc>=64 and cc<67) then grbp<="110";
	end if;
	if (cc=215 and ll=153) then grbp<="110";
	end if;
	if (cc=229 and ll=153) then grbp<="110";
	end if;
	if (cc=231 and ll=153) then grbp<="110";
	end if;
	if (cc=234 and ll=153) then grbp<="110";
	end if;
	if (cc=236 and ll=153) then grbp<="110";
	end if;
	if (cc=239 and ll=153) then grbp<="110";
	end if;
	if (ll=153 and cc>=239 and cc<246) then grbp<="110";
	end if;
	if (ll=153 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=154 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=141 and ll=154) then grbp<="110";
	end if;
	if (cc=220 and ll=154) then grbp<="110";
	end if;
	if (cc=223 and ll=154) then grbp<="110";
	end if;
	if (cc=240 and ll=154) then grbp<="110";
	end if;
	if (ll=154 and cc>=240 and cc<251) then grbp<="110";
	end if;
	if (ll=155 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=63 and ll=155) then grbp<="110";
	end if;
	if (cc=65 and ll=155) then grbp<="110";
	end if;
	if (cc=70 and ll=155) then grbp<="110";
	end if;
	if (cc=140 and ll=155) then grbp<="110";
	end if;
	if (cc=175 and ll=155) then grbp<="110";
	end if;
	if (cc=193 and ll=155) then grbp<="110";
	end if;
	if (cc=235 and ll=155) then grbp<="110";
	end if;
	if (cc=237 and ll=155) then grbp<="110";
	end if;
	if (cc=239 and ll=155) then grbp<="110";
	end if;
	if (cc=241 and ll=155) then grbp<="110";
	end if;
	if (ll=155 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=156 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=64 and ll=156) then grbp<="110";
	end if;
	if (ll=156 and cc>=64 and cc<66) then grbp<="110";
	end if;
	if (cc=187 and ll=156) then grbp<="110";
	end if;
	if (ll=156 and cc>=187 and cc<189) then grbp<="110";
	end if;
	if (cc=230 and ll=156) then grbp<="110";
	end if;
	if (cc=232 and ll=156) then grbp<="110";
	end if;
	if (ll=156 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (cc=241 and ll=156) then grbp<="110";
	end if;
	if (ll=156 and cc>=241 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=157) then grbp<="110";
	end if;
	if (ll=157 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=64 and ll=157) then grbp<="110";
	end if;
	if (ll=157 and cc>=64 and cc<66) then grbp<="110";
	end if;
	if (ll=157 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=218 and ll=157) then grbp<="110";
	end if;
	if (cc=237 and ll=157) then grbp<="110";
	end if;
	if (ll=157 and cc>=237 and cc<240) then grbp<="110";
	end if;
	if (ll=157 and cc>=241 and cc<245) then grbp<="110";
	end if;
	if (ll=157 and cc>=246 and cc<248) then grbp<="110";
	end if;
	if (ll=157 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=158 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=158) then grbp<="110";
	end if;
	if (cc=63 and ll=158) then grbp<="110";
	end if;
	if (cc=65 and ll=158) then grbp<="110";
	end if;
	if (ll=158 and cc>=65 and cc<67) then grbp<="110";
	end if;
	if (cc=138 and ll=158) then grbp<="110";
	end if;
	if (cc=184 and ll=158) then grbp<="110";
	end if;
	if (ll=158 and cc>=184 and cc<188) then grbp<="110";
	end if;
	if (cc=230 and ll=158) then grbp<="110";
	end if;
	if (ll=158 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (cc=239 and ll=158) then grbp<="110";
	end if;
	if (ll=158 and cc>=239 and cc<250) then grbp<="110";
	end if;
	if (ll=159 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=65 and ll=159) then grbp<="110";
	end if;
	if (ll=159 and cc>=65 and cc<67) then grbp<="110";
	end if;
	if (cc=182 and ll=159) then grbp<="110";
	end if;
	if (ll=159 and cc>=182 and cc<185) then grbp<="110";
	end if;
	if (ll=159 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=219 and ll=159) then grbp<="110";
	end if;
	if (cc=239 and ll=159) then grbp<="110";
	end if;
	if (cc=241 and ll=159) then grbp<="110";
	end if;
	if (cc=243 and ll=159) then grbp<="110";
	end if;
	if (ll=159 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=160 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=64 and ll=160) then grbp<="110";
	end if;
	if (cc=66 and ll=160) then grbp<="110";
	end if;
	if (ll=160 and cc>=66 and cc<68) then grbp<="110";
	end if;
	if (ll=160 and cc>=180 and cc<187) then grbp<="110";
	end if;
	if (ll=160 and cc>=217 and cc<219) then grbp<="110";
	end if;
	if (cc=222 and ll=160) then grbp<="110";
	end if;
	if (cc=235 and ll=160) then grbp<="110";
	end if;
	if (cc=237 and ll=160) then grbp<="110";
	end if;
	if (ll=160 and cc>=237 and cc<240) then grbp<="110";
	end if;
	if (ll=160 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (cc=249 and ll=160) then grbp<="110";
	end if;
	if (ll=160 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=161 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=161 and cc>=65 and cc<69) then grbp<="110";
	end if;
	if (cc=168 and ll=161) then grbp<="110";
	end if;
	if (cc=178 and ll=161) then grbp<="110";
	end if;
	if (ll=161 and cc>=178 and cc<184) then grbp<="110";
	end if;
	if (cc=230 and ll=161) then grbp<="110";
	end if;
	if (cc=235 and ll=161) then grbp<="110";
	end if;
	if (cc=240 and ll=161) then grbp<="110";
	end if;
	if (ll=161 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (cc=245 and ll=161) then grbp<="110";
	end if;
	if (ll=161 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=162 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=65 and ll=162) then grbp<="110";
	end if;
	if (cc=67 and ll=162) then grbp<="110";
	end if;
	if (ll=162 and cc>=67 and cc<69) then grbp<="110";
	end if;
	if (cc=178 and ll=162) then grbp<="110";
	end if;
	if (ll=162 and cc>=178 and cc<185) then grbp<="110";
	end if;
	if (cc=241 and ll=162) then grbp<="110";
	end if;
	if (ll=162 and cc>=241 and cc<243) then grbp<="110";
	end if;
	if (ll=162 and cc>=244 and cc<247) then grbp<="110";
	end if;
	if (ll=162 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=163 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=62 and ll=163) then grbp<="110";
	end if;
	if (cc=64 and ll=163) then grbp<="110";
	end if;
	if (cc=66 and ll=163) then grbp<="110";
	end if;
	if (ll=163 and cc>=66 and cc<70) then grbp<="110";
	end if;
	if (cc=134 and ll=163) then grbp<="110";
	end if;
	if (cc=166 and ll=163) then grbp<="110";
	end if;
	if (cc=178 and ll=163) then grbp<="110";
	end if;
	if (ll=163 and cc>=178 and cc<185) then grbp<="110";
	end if;
	if (ll=163 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (cc=240 and ll=163) then grbp<="110";
	end if;
	if (cc=244 and ll=163) then grbp<="110";
	end if;
	if (cc=246 and ll=163) then grbp<="110";
	end if;
	if (ll=163 and cc>=246 and cc<251) then grbp<="110";
	end if;
	if (ll=164 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=66 and ll=164) then grbp<="110";
	end if;
	if (ll=164 and cc>=66 and cc<68) then grbp<="110";
	end if;
	if (cc=71 and ll=164) then grbp<="110";
	end if;
	if (cc=165 and ll=164) then grbp<="110";
	end if;
	if (cc=178 and ll=164) then grbp<="110";
	end if;
	if (ll=164 and cc>=178 and cc<184) then grbp<="110";
	end if;
	if (cc=218 and ll=164) then grbp<="110";
	end if;
	if (cc=222 and ll=164) then grbp<="110";
	end if;
	if (cc=225 and ll=164) then grbp<="110";
	end if;
	if (cc=230 and ll=164) then grbp<="110";
	end if;
	if (ll=164 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=164 and cc>=239 and cc<243) then grbp<="110";
	end if;
	if (ll=164 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=165 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=165 and cc>=65 and cc<68) then grbp<="110";
	end if;
	if (cc=180 and ll=165) then grbp<="110";
	end if;
	if (ll=165 and cc>=180 and cc<182) then grbp<="110";
	end if;
	if (cc=216 and ll=165) then grbp<="110";
	end if;
	if (cc=222 and ll=165) then grbp<="110";
	end if;
	if (cc=225 and ll=165) then grbp<="110";
	end if;
	if (cc=229 and ll=165) then grbp<="110";
	end if;
	if (ll=165 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (cc=238 and ll=165) then grbp<="110";
	end if;
	if (cc=241 and ll=165) then grbp<="110";
	end if;
	if (cc=244 and ll=165) then grbp<="110";
	end if;
	if (ll=165 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (ll=165 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=166 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=65 and ll=166) then grbp<="110";
	end if;
	if (ll=166 and cc>=65 and cc<71) then grbp<="110";
	end if;
	if (ll=166 and cc>=179 and cc<183) then grbp<="110";
	end if;
	if (cc=233 and ll=166) then grbp<="110";
	end if;
	if (ll=166 and cc>=233 and cc<235) then grbp<="110";
	end if;
	if (ll=166 and cc>=239 and cc<242) then grbp<="110";
	end if;
	if (ll=166 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (ll=166 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=167 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=64 and ll=167) then grbp<="110";
	end if;
	if (cc=66 and ll=167) then grbp<="110";
	end if;
	if (ll=167 and cc>=66 and cc<69) then grbp<="110";
	end if;
	if (cc=179 and ll=167) then grbp<="110";
	end if;
	if (ll=167 and cc>=179 and cc<182) then grbp<="110";
	end if;
	if (cc=220 and ll=167) then grbp<="110";
	end if;
	if (cc=222 and ll=167) then grbp<="110";
	end if;
	if (cc=230 and ll=167) then grbp<="110";
	end if;
	if (ll=167 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (cc=243 and ll=167) then grbp<="110";
	end if;
	if (cc=245 and ll=167) then grbp<="110";
	end if;
	if (cc=247 and ll=167) then grbp<="110";
	end if;
	if (ll=167 and cc>=247 and cc<250) then grbp<="110";
	end if;
	if (ll=168 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=168 and cc>=67 and cc<71) then grbp<="110";
	end if;
	if (ll=168 and cc>=179 and cc<181) then grbp<="110";
	end if;
	if (cc=221 and ll=168) then grbp<="110";
	end if;
	if (cc=224 and ll=168) then grbp<="110";
	end if;
	if (cc=230 and ll=168) then grbp<="110";
	end if;
	if (cc=239 and ll=168) then grbp<="110";
	end if;
	if (ll=168 and cc>=239 and cc<242) then grbp<="110";
	end if;
	if (ll=168 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (ll=168 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=169 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=67 and ll=169) then grbp<="110";
	end if;
	if (ll=169 and cc>=67 and cc<71) then grbp<="110";
	end if;
	if (cc=184 and ll=169) then grbp<="110";
	end if;
	if (cc=219 and ll=169) then grbp<="110";
	end if;
	if (cc=224 and ll=169) then grbp<="110";
	end if;
	if (cc=230 and ll=169) then grbp<="110";
	end if;
	if (cc=239 and ll=169) then grbp<="110";
	end if;
	if (ll=169 and cc>=239 and cc<242) then grbp<="110";
	end if;
	if (ll=169 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=170 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (ll=170 and cc>=68 and cc<71) then grbp<="110";
	end if;
	if (ll=170 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (cc=227 and ll=170) then grbp<="110";
	end if;
	if (cc=232 and ll=170) then grbp<="110";
	end if;
	if (cc=240 and ll=170) then grbp<="110";
	end if;
	if (ll=170 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (ll=170 and cc>=244 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=171) then grbp<="110";
	end if;
	if (ll=171 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=171 and cc>=68 and cc<70) then grbp<="110";
	end if;
	if (cc=221 and ll=171) then grbp<="110";
	end if;
	if (ll=171 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (cc=229 and ll=171) then grbp<="110";
	end if;
	if (cc=237 and ll=171) then grbp<="110";
	end if;
	if (cc=240 and ll=171) then grbp<="110";
	end if;
	if (ll=171 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (cc=246 and ll=171) then grbp<="110";
	end if;
	if (ll=171 and cc>=246 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=172) then grbp<="110";
	end if;
	if (ll=172 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=68 and ll=172) then grbp<="110";
	end if;
	if (cc=236 and ll=172) then grbp<="110";
	end if;
	if (cc=242 and ll=172) then grbp<="110";
	end if;
	if (cc=244 and ll=172) then grbp<="110";
	end if;
	if (cc=246 and ll=172) then grbp<="110";
	end if;
	if (ll=172 and cc>=246 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=173) then grbp<="110";
	end if;
	if (ll=173 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=180 and ll=173) then grbp<="110";
	end if;
	if (cc=214 and ll=173) then grbp<="110";
	end if;
	if (cc=220 and ll=173) then grbp<="110";
	end if;
	if (cc=222 and ll=173) then grbp<="110";
	end if;
	if (cc=236 and ll=173) then grbp<="110";
	end if;
	if (cc=238 and ll=173) then grbp<="110";
	end if;
	if (cc=242 and ll=173) then grbp<="110";
	end if;
	if (ll=173 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (cc=248 and ll=173) then grbp<="110";
	end if;
	if (ll=173 and cc>=248 and cc<251) then grbp<="110";
	end if;
	if (ll=174 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=179 and ll=174) then grbp<="110";
	end if;
	if (cc=217 and ll=174) then grbp<="110";
	end if;
	if (cc=225 and ll=174) then grbp<="110";
	end if;
	if (cc=229 and ll=174) then grbp<="110";
	end if;
	if (ll=174 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (cc=235 and ll=174) then grbp<="110";
	end if;
	if (ll=174 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (cc=246 and ll=174) then grbp<="110";
	end if;
	if (ll=174 and cc>=246 and cc<250) then grbp<="110";
	end if;
	if (ll=175 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=224 and ll=175) then grbp<="110";
	end if;
	if (cc=226 and ll=175) then grbp<="110";
	end if;
	if (cc=228 and ll=175) then grbp<="110";
	end if;
	if (cc=235 and ll=175) then grbp<="110";
	end if;
	if (cc=241 and ll=175) then grbp<="110";
	end if;
	if (cc=244 and ll=175) then grbp<="110";
	end if;
	if (ll=175 and cc>=244 and cc<250) then grbp<="110";
	end if;
	if (ll=176 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=176 and cc>=69 and cc<71) then grbp<="110";
	end if;
	if (cc=218 and ll=176) then grbp<="110";
	end if;
	if (cc=220 and ll=176) then grbp<="110";
	end if;
	if (cc=225 and ll=176) then grbp<="110";
	end if;
	if (cc=229 and ll=176) then grbp<="110";
	end if;
	if (cc=235 and ll=176) then grbp<="110";
	end if;
	if (ll=176 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (ll=176 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=176 and cc>=243 and cc<251) then grbp<="110";
	end if;
	if (ll=177 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=220 and ll=177) then grbp<="110";
	end if;
	if (cc=228 and ll=177) then grbp<="110";
	end if;
	if (cc=238 and ll=177) then grbp<="110";
	end if;
	if (ll=177 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=177 and cc>=242 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=178) then grbp<="110";
	end if;
	if (ll=178 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=222 and ll=178) then grbp<="110";
	end if;
	if (cc=228 and ll=178) then grbp<="110";
	end if;
	if (cc=238 and ll=178) then grbp<="110";
	end if;
	if (ll=178 and cc>=238 and cc<251) then grbp<="110";
	end if;
	if (ll=179 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=213 and ll=179) then grbp<="110";
	end if;
	if (ll=179 and cc>=213 and cc<217) then grbp<="110";
	end if;
	if (ll=179 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=179 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (cc=233 and ll=179) then grbp<="110";
	end if;
	if (cc=240 and ll=179) then grbp<="110";
	end if;
	if (cc=243 and ll=179) then grbp<="110";
	end if;
	if (cc=245 and ll=179) then grbp<="110";
	end if;
	if (ll=179 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (cc=250 and ll=179) then grbp<="110";
	end if;
	if (cc=17 and ll=180) then grbp<="110";
	end if;
	if (ll=180 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=180 and cc>=68 and cc<70) then grbp<="110";
	end if;
	if (ll=180 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=222 and ll=180) then grbp<="110";
	end if;
	if (ll=180 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=180 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=180 and cc>=231 and cc<234) then grbp<="110";
	end if;
	if (ll=180 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (cc=243 and ll=180) then grbp<="110";
	end if;
	if (ll=180 and cc>=243 and cc<246) then grbp<="110";
	end if;
	if (ll=180 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=181 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=215 and ll=181) then grbp<="110";
	end if;
	if (cc=217 and ll=181) then grbp<="110";
	end if;
	if (cc=224 and ll=181) then grbp<="110";
	end if;
	if (cc=226 and ll=181) then grbp<="110";
	end if;
	if (cc=233 and ll=181) then grbp<="110";
	end if;
	if (cc=239 and ll=181) then grbp<="110";
	end if;
	if (cc=241 and ll=181) then grbp<="110";
	end if;
	if (cc=243 and ll=181) then grbp<="110";
	end if;
	if (cc=245 and ll=181) then grbp<="110";
	end if;
	if (cc=247 and ll=181) then grbp<="110";
	end if;
	if (ll=181 and cc>=247 and cc<250) then grbp<="110";
	end if;
	if (ll=182 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=166 and ll=182) then grbp<="110";
	end if;
	if (cc=212 and ll=182) then grbp<="110";
	end if;
	if (ll=182 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (ll=182 and cc>=215 and cc<217) then grbp<="110";
	end if;
	if (cc=225 and ll=182) then grbp<="110";
	end if;
	if (ll=182 and cc>=225 and cc<229) then grbp<="110";
	end if;
	if (cc=242 and ll=182) then grbp<="110";
	end if;
	if (cc=244 and ll=182) then grbp<="110";
	end if;
	if (ll=182 and cc>=244 and cc<250) then grbp<="110";
	end if;
	if (ll=183 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=68 and ll=183) then grbp<="110";
	end if;
	if (cc=212 and ll=183) then grbp<="110";
	end if;
	if (ll=183 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=218 and ll=183) then grbp<="110";
	end if;
	if (cc=225 and ll=183) then grbp<="110";
	end if;
	if (ll=183 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (cc=236 and ll=183) then grbp<="110";
	end if;
	if (cc=240 and ll=183) then grbp<="110";
	end if;
	if (ll=183 and cc>=240 and cc<245) then grbp<="110";
	end if;
	if (ll=183 and cc>=246 and cc<250) then grbp<="110";
	end if;
	if (ll=184 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=121 and ll=184) then grbp<="110";
	end if;
	if (cc=211 and ll=184) then grbp<="110";
	end if;
	if (ll=184 and cc>=211 and cc<215) then grbp<="110";
	end if;
	if (ll=184 and cc>=216 and cc<218) then grbp<="110";
	end if;
	if (cc=225 and ll=184) then grbp<="110";
	end if;
	if (ll=184 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (cc=231 and ll=184) then grbp<="110";
	end if;
	if (ll=184 and cc>=231 and cc<234) then grbp<="110";
	end if;
	if (cc=240 and ll=184) then grbp<="110";
	end if;
	if (cc=242 and ll=184) then grbp<="110";
	end if;
	if (ll=184 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (ll=184 and cc>=246 and cc<250) then grbp<="110";
	end if;
	if (ll=185 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=212 and ll=185) then grbp<="110";
	end if;
	if (ll=185 and cc>=212 and cc<216) then grbp<="110";
	end if;
	if (cc=220 and ll=185) then grbp<="110";
	end if;
	if (ll=185 and cc>=220 and cc<224) then grbp<="110";
	end if;
	if (ll=185 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=185 and cc>=229 and cc<233) then grbp<="110";
	end if;
	if (cc=242 and ll=185) then grbp<="110";
	end if;
	if (ll=185 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (ll=185 and cc>=246 and cc<250) then grbp<="110";
	end if;
	if (ll=186 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=212 and ll=186) then grbp<="110";
	end if;
	if (cc=215 and ll=186) then grbp<="110";
	end if;
	if (cc=220 and ll=186) then grbp<="110";
	end if;
	if (ll=186 and cc>=220 and cc<223) then grbp<="110";
	end if;
	if (ll=186 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (cc=238 and ll=186) then grbp<="110";
	end if;
	if (ll=186 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=186 and cc>=241 and cc<251) then grbp<="110";
	end if;
	if (ll=187 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=119 and ll=187) then grbp<="110";
	end if;
	if (cc=210 and ll=187) then grbp<="110";
	end if;
	if (cc=212 and ll=187) then grbp<="110";
	end if;
	if (ll=187 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (ll=187 and cc>=215 and cc<223) then grbp<="110";
	end if;
	if (ll=187 and cc>=225 and cc<229) then grbp<="110";
	end if;
	if (cc=238 and ll=187) then grbp<="110";
	end if;
	if (ll=187 and cc>=238 and cc<245) then grbp<="110";
	end if;
	if (ll=187 and cc>=246 and cc<250) then grbp<="110";
	end if;
	if (ll=188 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=65 and ll=188) then grbp<="110";
	end if;
	if (cc=141 and ll=188) then grbp<="110";
	end if;
	if (cc=167 and ll=188) then grbp<="110";
	end if;
	if (cc=212 and ll=188) then grbp<="110";
	end if;
	if (ll=188 and cc>=212 and cc<219) then grbp<="110";
	end if;
	if (cc=223 and ll=188) then grbp<="110";
	end if;
	if (ll=188 and cc>=223 and cc<228) then grbp<="110";
	end if;
	if (cc=240 and ll=188) then grbp<="110";
	end if;
	if (ll=188 and cc>=240 and cc<245) then grbp<="110";
	end if;
	if (cc=248 and ll=188) then grbp<="110";
	end if;
	if (cc=17 and ll=189) then grbp<="110";
	end if;
	if (ll=189 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=118 and ll=189) then grbp<="110";
	end if;
	if (cc=167 and ll=189) then grbp<="110";
	end if;
	if (cc=212 and ll=189) then grbp<="110";
	end if;
	if (cc=214 and ll=189) then grbp<="110";
	end if;
	if (ll=189 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=189 and cc>=217 and cc<221) then grbp<="110";
	end if;
	if (ll=189 and cc>=222 and cc<232) then grbp<="110";
	end if;
	if (cc=238 and ll=189) then grbp<="110";
	end if;
	if (cc=241 and ll=189) then grbp<="110";
	end if;
	if (ll=189 and cc>=241 and cc<243) then grbp<="110";
	end if;
	if (ll=189 and cc>=244 and cc<249) then grbp<="110";
	end if;
	if (ll=190 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=212 and ll=190) then grbp<="110";
	end if;
	if (ll=190 and cc>=212 and cc<215) then grbp<="110";
	end if;
	if (ll=190 and cc>=220 and cc<223) then grbp<="110";
	end if;
	if (cc=228 and ll=190) then grbp<="110";
	end if;
	if (ll=190 and cc>=228 and cc<232) then grbp<="110";
	end if;
	if (cc=241 and ll=190) then grbp<="110";
	end if;
	if (ll=190 and cc>=241 and cc<250) then grbp<="110";
	end if;
	if (ll=191 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=139 and ll=191) then grbp<="110";
	end if;
	if (cc=141 and ll=191) then grbp<="110";
	end if;
	if (cc=209 and ll=191) then grbp<="110";
	end if;
	if (cc=214 and ll=191) then grbp<="110";
	end if;
	if (ll=191 and cc>=214 and cc<221) then grbp<="110";
	end if;
	if (ll=191 and cc>=224 and cc<228) then grbp<="110";
	end if;
	if (cc=231 and ll=191) then grbp<="110";
	end if;
	if (ll=191 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (cc=238 and ll=191) then grbp<="110";
	end if;
	if (ll=191 and cc>=238 and cc<241) then grbp<="110";
	end if;
	if (ll=191 and cc>=242 and cc<248) then grbp<="110";
	end if;
	if (cc=17 and ll=192) then grbp<="110";
	end if;
	if (ll=192 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=209 and ll=192) then grbp<="110";
	end if;
	if (ll=192 and cc>=209 and cc<211) then grbp<="110";
	end if;
	if (cc=214 and ll=192) then grbp<="110";
	end if;
	if (ll=192 and cc>=214 and cc<222) then grbp<="110";
	end if;
	if (ll=192 and cc>=223 and cc<227) then grbp<="110";
	end if;
	if (ll=192 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (cc=234 and ll=192) then grbp<="110";
	end if;
	if (cc=236 and ll=192) then grbp<="110";
	end if;
	if (cc=239 and ll=192) then grbp<="110";
	end if;
	if (cc=241 and ll=192) then grbp<="110";
	end if;
	if (cc=243 and ll=192) then grbp<="110";
	end if;
	if (ll=192 and cc>=243 and cc<246) then grbp<="110";
	end if;
	if (ll=192 and cc>=247 and cc<250) then grbp<="110";
	end if;
	if (ll=193 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=116 and ll=193) then grbp<="110";
	end if;
	if (cc=140 and ll=193) then grbp<="110";
	end if;
	if (cc=209 and ll=193) then grbp<="110";
	end if;
	if (cc=214 and ll=193) then grbp<="110";
	end if;
	if (ll=193 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=193 and cc>=217 and cc<222) then grbp<="110";
	end if;
	if (ll=193 and cc>=223 and cc<226) then grbp<="110";
	end if;
	if (cc=233 and ll=193) then grbp<="110";
	end if;
	if (ll=193 and cc>=233 and cc<237) then grbp<="110";
	end if;
	if (ll=193 and cc>=239 and cc<246) then grbp<="110";
	end if;
	if (ll=193 and cc>=247 and cc<250) then grbp<="110";
	end if;
	if (ll=194 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=120 and ll=194) then grbp<="110";
	end if;
	if (cc=138 and ll=194) then grbp<="110";
	end if;
	if (ll=194 and cc>=138 and cc<140) then grbp<="110";
	end if;
	if (ll=194 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=217 and ll=194) then grbp<="110";
	end if;
	if (cc=224 and ll=194) then grbp<="110";
	end if;
	if (cc=226 and ll=194) then grbp<="110";
	end if;
	if (ll=194 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (cc=231 and ll=194) then grbp<="110";
	end if;
	if (cc=233 and ll=194) then grbp<="110";
	end if;
	if (cc=235 and ll=194) then grbp<="110";
	end if;
	if (ll=194 and cc>=235 and cc<238) then grbp<="110";
	end if;
	if (ll=194 and cc>=239 and cc<250) then grbp<="110";
	end if;
	if (ll=195 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=195 and cc>=23 and cc<28) then grbp<="110";
	end if;
	if (cc=115 and ll=195) then grbp<="110";
	end if;
	if (cc=213 and ll=195) then grbp<="110";
	end if;
	if (cc=215 and ll=195) then grbp<="110";
	end if;
	if (cc=217 and ll=195) then grbp<="110";
	end if;
	if (cc=220 and ll=195) then grbp<="110";
	end if;
	if (cc=222 and ll=195) then grbp<="110";
	end if;
	if (ll=195 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=195 and cc>=225 and cc<228) then grbp<="110";
	end if;
	if (ll=195 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (cc=235 and ll=195) then grbp<="110";
	end if;
	if (cc=238 and ll=195) then grbp<="110";
	end if;
	if (ll=195 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (cc=246 and ll=195) then grbp<="110";
	end if;
	if (ll=195 and cc>=246 and cc<249) then grbp<="110";
	end if;
	if (ll=196 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=119 and ll=196) then grbp<="110";
	end if;
	if (ll=196 and cc>=119 and cc<121) then grbp<="110";
	end if;
	if (cc=210 and ll=196) then grbp<="110";
	end if;
	if (cc=217 and ll=196) then grbp<="110";
	end if;
	if (cc=220 and ll=196) then grbp<="110";
	end if;
	if (cc=223 and ll=196) then grbp<="110";
	end if;
	if (cc=225 and ll=196) then grbp<="110";
	end if;
	if (ll=196 and cc>=225 and cc<229) then grbp<="110";
	end if;
	if (ll=196 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (ll=196 and cc>=241 and cc<250) then grbp<="110";
	end if;
	if (ll=197 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=197 and cc>=119 and cc<121) then grbp<="110";
	end if;
	if (cc=208 and ll=197) then grbp<="110";
	end if;
	if (cc=210 and ll=197) then grbp<="110";
	end if;
	if (cc=212 and ll=197) then grbp<="110";
	end if;
	if (cc=215 and ll=197) then grbp<="110";
	end if;
	if (ll=197 and cc>=215 and cc<218) then grbp<="110";
	end if;
	if (cc=224 and ll=197) then grbp<="110";
	end if;
	if (ll=197 and cc>=224 and cc<228) then grbp<="110";
	end if;
	if (cc=231 and ll=197) then grbp<="110";
	end if;
	if (ll=197 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (ll=197 and cc>=242 and cc<244) then grbp<="110";
	end if;
	if (ll=197 and cc>=245 and cc<249) then grbp<="110";
	end if;
	if (cc=17 and ll=198) then grbp<="110";
	end if;
	if (ll=198 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=198 and cc>=118 and cc<120) then grbp<="110";
	end if;
	if (cc=216 and ll=198) then grbp<="110";
	end if;
	if (cc=218 and ll=198) then grbp<="110";
	end if;
	if (cc=223 and ll=198) then grbp<="110";
	end if;
	if (ll=198 and cc>=223 and cc<227) then grbp<="110";
	end if;
	if (cc=230 and ll=198) then grbp<="110";
	end if;
	if (ll=198 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (cc=235 and ll=198) then grbp<="110";
	end if;
	if (cc=245 and ll=198) then grbp<="110";
	end if;
	if (ll=198 and cc>=245 and cc<251) then grbp<="110";
	end if;
	if (ll=199 and cc>=16 and cc<28) then grbp<="110";
	end if;
	if (cc=208 and ll=199) then grbp<="110";
	end if;
	if (ll=199 and cc>=208 and cc<210) then grbp<="110";
	end if;
	if (cc=216 and ll=199) then grbp<="110";
	end if;
	if (ll=199 and cc>=216 and cc<219) then grbp<="110";
	end if;
	if (ll=199 and cc>=226 and cc<234) then grbp<="110";
	end if;
	if (ll=199 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (ll=199 and cc>=247 and cc<251) then grbp<="110";
	end if;
	if (ll=200 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=200 and cc>=24 and cc<28) then grbp<="110";
	end if;
	if (cc=117 and ll=200) then grbp<="110";
	end if;
	if (cc=209 and ll=200) then grbp<="110";
	end if;
	if (ll=200 and cc>=209 and cc<212) then grbp<="110";
	end if;
	if (cc=216 and ll=200) then grbp<="110";
	end if;
	if (ll=200 and cc>=216 and cc<219) then grbp<="110";
	end if;
	if (ll=200 and cc>=226 and cc<232) then grbp<="110";
	end if;
	if (cc=249 and ll=200) then grbp<="110";
	end if;
	if (ll=200 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=201 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=68 and ll=201) then grbp<="110";
	end if;
	if (ll=201 and cc>=68 and cc<70) then grbp<="110";
	end if;
	if (cc=209 and ll=201) then grbp<="110";
	end if;
	if (cc=213 and ll=201) then grbp<="110";
	end if;
	if (ll=201 and cc>=213 and cc<219) then grbp<="110";
	end if;
	if (cc=227 and ll=201) then grbp<="110";
	end if;
	if (ll=201 and cc>=227 and cc<234) then grbp<="110";
	end if;
	if (ll=202 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=121 and ll=202) then grbp<="110";
	end if;
	if (cc=207 and ll=202) then grbp<="110";
	end if;
	if (ll=202 and cc>=207 and cc<209) then grbp<="110";
	end if;
	if (cc=212 and ll=202) then grbp<="110";
	end if;
	if (cc=215 and ll=202) then grbp<="110";
	end if;
	if (ll=202 and cc>=215 and cc<220) then grbp<="110";
	end if;
	if (cc=227 and ll=202) then grbp<="110";
	end if;
	if (ll=202 and cc>=227 and cc<235) then grbp<="110";
	end if;
	if (ll=203 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=203 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=207 and ll=203) then grbp<="110";
	end if;
	if (ll=203 and cc>=207 and cc<211) then grbp<="110";
	end if;
	if (ll=203 and cc>=213 and cc<221) then grbp<="110";
	end if;
	if (ll=203 and cc>=226 and cc<231) then grbp<="110";
	end if;
	if (ll=203 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (cc=237 and ll=203) then grbp<="110";
	end if;
	if (ll=203 and cc>=237 and cc<239) then grbp<="110";
	end if;
	if (ll=204 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=115 and ll=204) then grbp<="110";
	end if;
	if (cc=120 and ll=204) then grbp<="110";
	end if;
	if (cc=207 and ll=204) then grbp<="110";
	end if;
	if (cc=209 and ll=204) then grbp<="110";
	end if;
	if (cc=211 and ll=204) then grbp<="110";
	end if;
	if (ll=204 and cc>=211 and cc<214) then grbp<="110";
	end if;
	if (ll=204 and cc>=215 and cc<222) then grbp<="110";
	end if;
	if (ll=204 and cc>=223 and cc<231) then grbp<="110";
	end if;
	if (ll=204 and cc>=232 and cc<237) then grbp<="110";
	end if;
	if (ll=205 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=206 and ll=205) then grbp<="110";
	end if;
	if (ll=205 and cc>=206 and cc<212) then grbp<="110";
	end if;
	if (ll=205 and cc>=213 and cc<217) then grbp<="110";
	end if;
	if (ll=205 and cc>=218 and cc<221) then grbp<="110";
	end if;
	if (ll=205 and cc>=223 and cc<233) then grbp<="110";
	end if;
	if (ll=205 and cc>=234 and cc<236) then grbp<="110";
	end if;
	if (cc=17 and ll=206) then grbp<="110";
	end if;
	if (ll=206 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=206 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (ll=206 and cc>=71 and cc<73) then grbp<="110";
	end if;
	if (cc=114 and ll=206) then grbp<="110";
	end if;
	if (cc=206 and ll=206) then grbp<="110";
	end if;
	if (ll=206 and cc>=206 and cc<215) then grbp<="110";
	end if;
	if (ll=206 and cc>=216 and cc<219) then grbp<="110";
	end if;
	if (cc=226 and ll=206) then grbp<="110";
	end if;
	if (ll=206 and cc>=226 and cc<235) then grbp<="110";
	end if;
	if (ll=207 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=207 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (cc=163 and ll=207) then grbp<="110";
	end if;
	if (cc=206 and ll=207) then grbp<="110";
	end if;
	if (ll=207 and cc>=206 and cc<214) then grbp<="110";
	end if;
	if (ll=207 and cc>=216 and cc<223) then grbp<="110";
	end if;
	if (ll=207 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (ll=207 and cc>=227 and cc<234) then grbp<="110";
	end if;
	if (cc=17 and ll=208) then grbp<="110";
	end if;
	if (ll=208 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=114 and ll=208) then grbp<="110";
	end if;
	if (cc=125 and ll=208) then grbp<="110";
	end if;
	if (cc=132 and ll=208) then grbp<="110";
	end if;
	if (cc=144 and ll=208) then grbp<="110";
	end if;
	if (cc=162 and ll=208) then grbp<="110";
	end if;
	if (cc=206 and ll=208) then grbp<="110";
	end if;
	if (ll=208 and cc>=206 and cc<211) then grbp<="110";
	end if;
	if (ll=208 and cc>=212 and cc<215) then grbp<="110";
	end if;
	if (cc=218 and ll=208) then grbp<="110";
	end if;
	if (ll=208 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=208 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=208 and cc>=224 and cc<231) then grbp<="110";
	end if;
	if (ll=208 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (cc=242 and ll=208) then grbp<="110";
	end if;
	if (cc=18 and ll=209) then grbp<="110";
	end if;
	if (ll=209 and cc>=18 and cc<28) then grbp<="110";
	end if;
	if (cc=109 and ll=209) then grbp<="110";
	end if;
	if (cc=113 and ll=209) then grbp<="110";
	end if;
	if (cc=119 and ll=209) then grbp<="110";
	end if;
	if (cc=161 and ll=209) then grbp<="110";
	end if;
	if (cc=206 and ll=209) then grbp<="110";
	end if;
	if (ll=209 and cc>=206 and cc<209) then grbp<="110";
	end if;
	if (cc=212 and ll=209) then grbp<="110";
	end if;
	if (cc=214 and ll=209) then grbp<="110";
	end if;
	if (ll=209 and cc>=214 and cc<223) then grbp<="110";
	end if;
	if (ll=209 and cc>=224 and cc<235) then grbp<="110";
	end if;
	if (cc=242 and ll=209) then grbp<="110";
	end if;
	if (cc=17 and ll=210) then grbp<="110";
	end if;
	if (ll=210 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=63 and ll=210) then grbp<="110";
	end if;
	if (cc=145 and ll=210) then grbp<="110";
	end if;
	if (cc=205 and ll=210) then grbp<="110";
	end if;
	if (ll=210 and cc>=205 and cc<234) then grbp<="110";
	end if;
	if (ll=210 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (cc=17 and ll=211) then grbp<="110";
	end if;
	if (ll=211 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=63 and ll=211) then grbp<="110";
	end if;
	if (ll=211 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=113 and ll=211) then grbp<="110";
	end if;
	if (cc=205 and ll=211) then grbp<="110";
	end if;
	if (ll=211 and cc>=205 and cc<209) then grbp<="110";
	end if;
	if (ll=211 and cc>=210 and cc<234) then grbp<="110";
	end if;
	if (ll=211 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (cc=245 and ll=211) then grbp<="110";
	end if;
	if (cc=17 and ll=212) then grbp<="110";
	end if;
	if (ll=212 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=212 and cc>=59 and cc<61) then grbp<="110";
	end if;
	if (ll=212 and cc>=63 and cc<66) then grbp<="110";
	end if;
	if (cc=149 and ll=212) then grbp<="110";
	end if;
	if (cc=205 and ll=212) then grbp<="110";
	end if;
	if (ll=212 and cc>=205 and cc<221) then grbp<="110";
	end if;
	if (ll=212 and cc>=222 and cc<238) then grbp<="110";
	end if;
	if (ll=212 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (ll=213 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=213 and cc>=59 and cc<62) then grbp<="110";
	end if;
	if (ll=213 and cc>=63 and cc<65) then grbp<="110";
	end if;
	if (cc=159 and ll=213) then grbp<="110";
	end if;
	if (cc=205 and ll=213) then grbp<="110";
	end if;
	if (cc=207 and ll=213) then grbp<="110";
	end if;
	if (cc=209 and ll=213) then grbp<="110";
	end if;
	if (ll=213 and cc>=209 and cc<231) then grbp<="110";
	end if;
	if (ll=213 and cc>=232 and cc<236) then grbp<="110";
	end if;
	if (ll=213 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (ll=214 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=149 and ll=214) then grbp<="110";
	end if;
	if (cc=205 and ll=214) then grbp<="110";
	end if;
	if (ll=214 and cc>=205 and cc<209) then grbp<="110";
	end if;
	if (ll=214 and cc>=210 and cc<235) then grbp<="110";
	end if;
	if (cc=238 and ll=214) then grbp<="110";
	end if;
	if (cc=242 and ll=214) then grbp<="110";
	end if;
	if (cc=17 and ll=215) then grbp<="110";
	end if;
	if (ll=215 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=215 and cc>=62 and cc<64) then grbp<="110";
	end if;
	if (cc=149 and ll=215) then grbp<="110";
	end if;
	if (cc=158 and ll=215) then grbp<="110";
	end if;
	if (cc=205 and ll=215) then grbp<="110";
	end if;
	if (ll=215 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (ll=215 and cc>=209 and cc<213) then grbp<="110";
	end if;
	if (ll=215 and cc>=214 and cc<234) then grbp<="110";
	end if;
	if (cc=237 and ll=215) then grbp<="110";
	end if;
	if (ll=215 and cc>=237 and cc<242) then grbp<="110";
	end if;
	if (ll=216 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=149 and ll=216) then grbp<="110";
	end if;
	if (cc=204 and ll=216) then grbp<="110";
	end if;
	if (ll=216 and cc>=204 and cc<233) then grbp<="110";
	end if;
	if (ll=216 and cc>=235 and cc<239) then grbp<="110";
	end if;
	if (cc=17 and ll=217) then grbp<="110";
	end if;
	if (ll=217 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=61 and ll=217) then grbp<="110";
	end if;
	if (cc=106 and ll=217) then grbp<="110";
	end if;
	if (cc=205 and ll=217) then grbp<="110";
	end if;
	if (ll=217 and cc>=205 and cc<235) then grbp<="110";
	end if;
	if (ll=217 and cc>=237 and cc<239) then grbp<="110";
	end if;
	if (ll=218 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=60 and ll=218) then grbp<="110";
	end if;
	if (cc=204 and ll=218) then grbp<="110";
	end if;
	if (ll=218 and cc>=204 and cc<234) then grbp<="110";
	end if;
	if (ll=218 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (ll=218 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=219 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=60 and ll=219) then grbp<="110";
	end if;
	if (cc=118 and ll=219) then grbp<="110";
	end if;
	if (cc=204 and ll=219) then grbp<="110";
	end if;
	if (ll=219 and cc>=204 and cc<234) then grbp<="110";
	end if;
	if (cc=237 and ll=219) then grbp<="110";
	end if;
	if (cc=17 and ll=220) then grbp<="110";
	end if;
	if (ll=220 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=220 and cc>=25 and cc<28) then grbp<="110";
	end if;
	if (cc=105 and ll=220) then grbp<="110";
	end if;
	if (cc=203 and ll=220) then grbp<="110";
	end if;
	if (ll=220 and cc>=203 and cc<233) then grbp<="110";
	end if;
	if (ll=220 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (ll=221 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (cc=155 and ll=221) then grbp<="110";
	end if;
	if (cc=203 and ll=221) then grbp<="110";
	end if;
	if (ll=221 and cc>=203 and cc<233) then grbp<="110";
	end if;
	if (cc=17 and ll=222) then grbp<="110";
	end if;
	if (ll=222 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=203 and ll=222) then grbp<="110";
	end if;
	if (cc=205 and ll=222) then grbp<="110";
	end if;
	if (ll=222 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (ll=222 and cc>=209 and cc<234) then grbp<="110";
	end if;
	if (cc=250 and ll=222) then grbp<="110";
	end if;
	if (cc=17 and ll=223) then grbp<="110";
	end if;
	if (ll=223 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=223 and cc>=26 and cc<28) then grbp<="110";
	end if;
	if (ll=223 and cc>=58 and cc<60) then grbp<="110";
	end if;
	if (cc=203 and ll=223) then grbp<="110";
	end if;
	if (ll=223 and cc>=203 and cc<208) then grbp<="110";
	end if;
	if (ll=223 and cc>=209 and cc<231) then grbp<="110";
	end if;
	if (cc=17 and ll=224) then grbp<="110";
	end if;
	if (ll=224 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=203 and ll=224) then grbp<="110";
	end if;
	if (ll=224 and cc>=203 and cc<212) then grbp<="110";
	end if;
	if (cc=215 and ll=224) then grbp<="110";
	end if;
	if (ll=224 and cc>=215 and cc<230) then grbp<="110";
	end if;
	if (cc=17 and ll=225) then grbp<="110";
	end if;
	if (ll=225 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=225 and cc>=25 and cc<28) then grbp<="110";
	end if;
	if (cc=115 and ll=225) then grbp<="110";
	end if;
	if (cc=137 and ll=225) then grbp<="110";
	end if;
	if (cc=149 and ll=225) then grbp<="110";
	end if;
	if (cc=202 and ll=225) then grbp<="110";
	end if;
	if (ll=225 and cc>=202 and cc<230) then grbp<="110";
	end if;
	if (ll=225 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (cc=17 and ll=226) then grbp<="110";
	end if;
	if (ll=226 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=226 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=202 and ll=226) then grbp<="110";
	end if;
	if (ll=226 and cc>=202 and cc<216) then grbp<="110";
	end if;
	if (ll=226 and cc>=217 and cc<227) then grbp<="110";
	end if;
	if (ll=226 and cc>=228 and cc<232) then grbp<="110";
	end if;
	if (cc=17 and ll=227) then grbp<="110";
	end if;
	if (ll=227 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=227 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=227 and cc>=204 and cc<216) then grbp<="110";
	end if;
	if (ll=227 and cc>=218 and cc<226) then grbp<="110";
	end if;
	if (cc=232 and ll=227) then grbp<="110";
	end if;
	if (cc=243 and ll=227) then grbp<="110";
	end if;
	if (cc=245 and ll=227) then grbp<="110";
	end if;
	if (cc=17 and ll=228) then grbp<="110";
	end if;
	if (ll=228 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (cc=26 and ll=228) then grbp<="110";
	end if;
	if (ll=228 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=204 and ll=228) then grbp<="110";
	end if;
	if (ll=228 and cc>=204 and cc<212) then grbp<="110";
	end if;
	if (ll=228 and cc>=213 and cc<216) then grbp<="110";
	end if;
	if (ll=228 and cc>=218 and cc<228) then grbp<="110";
	end if;
	if (ll=228 and cc>=243 and cc<245) then grbp<="110";
	end if;
	if (ll=229 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=229 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (cc=56 and ll=229) then grbp<="110";
	end if;
	if (cc=202 and ll=229) then grbp<="110";
	end if;
	if (cc=204 and ll=229) then grbp<="110";
	end if;
	if (ll=229 and cc>=204 and cc<210) then grbp<="110";
	end if;
	if (cc=215 and ll=229) then grbp<="110";
	end if;
	if (cc=218 and ll=229) then grbp<="110";
	end if;
	if (ll=229 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=229 and cc>=221 and cc<226) then grbp<="110";
	end if;
	if (cc=242 and ll=229) then grbp<="110";
	end if;
	if (cc=17 and ll=230) then grbp<="110";
	end if;
	if (ll=230 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=230 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=230 and cc>=202 and cc<211) then grbp<="110";
	end if;
	if (ll=230 and cc>=212 and cc<215) then grbp<="110";
	end if;
	if (ll=230 and cc>=216 and cc<226) then grbp<="110";
	end if;
	if (ll=230 and cc>=241 and cc<243) then grbp<="110";
	end if;
	if (ll=231 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=203 and ll=231) then grbp<="110";
	end if;
	if (ll=231 and cc>=203 and cc<226) then grbp<="110";
	end if;
	if (ll=231 and cc>=240 and cc<242) then grbp<="110";
	end if;
	if (cc=17 and ll=232) then grbp<="110";
	end if;
	if (ll=232 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=232 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=232 and cc>=201 and cc<224) then grbp<="110";
	end if;
	if (ll=232 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=232 and cc>=238 and cc<241) then grbp<="110";
	end if;
	if (cc=17 and ll=233) then grbp<="110";
	end if;
	if (ll=233 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=233 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=203 and ll=233) then grbp<="110";
	end if;
	if (ll=233 and cc>=203 and cc<210) then grbp<="110";
	end if;
	if (cc=213 and ll=233) then grbp<="110";
	end if;
	if (cc=215 and ll=233) then grbp<="110";
	end if;
	if (ll=233 and cc>=215 and cc<225) then grbp<="110";
	end if;
	if (ll=233 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=234 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=234 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=201 and ll=234) then grbp<="110";
	end if;
	if (ll=234 and cc>=201 and cc<206) then grbp<="110";
	end if;
	if (cc=209 and ll=234) then grbp<="110";
	end if;
	if (ll=234 and cc>=209 and cc<214) then grbp<="110";
	end if;
	if (cc=217 and ll=234) then grbp<="110";
	end if;
	if (ll=234 and cc>=217 and cc<224) then grbp<="110";
	end if;
	if (ll=235 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=235 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=201 and ll=235) then grbp<="110";
	end if;
	if (ll=235 and cc>=201 and cc<210) then grbp<="110";
	end if;
	if (ll=235 and cc>=211 and cc<224) then grbp<="110";
	end if;
	if (ll=236 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=236 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (ll=236 and cc>=201 and cc<223) then grbp<="110";
	end if;
	if (ll=237 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=237 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=237 and cc>=200 and cc<212) then grbp<="110";
	end if;
	if (ll=237 and cc>=213 and cc<217) then grbp<="110";
	end if;
	if (ll=237 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=238 and cc>=18 and cc<22) then grbp<="110";
	end if;
	if (cc=25 and ll=238) then grbp<="110";
	end if;
	if (ll=238 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=159 and ll=238) then grbp<="110";
	end if;
	if (cc=200 and ll=238) then grbp<="110";
	end if;
	if (cc=202 and ll=238) then grbp<="110";
	end if;
	if (ll=238 and cc>=202 and cc<209) then grbp<="110";
	end if;
	if (ll=238 and cc>=211 and cc<217) then grbp<="110";
	end if;
	if (ll=238 and cc>=218 and cc<222) then grbp<="110";
	end if;
	if (cc=17 and ll=239) then grbp<="110";
	end if;
	if (ll=239 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=239 and cc>=23 and cc<25) then grbp<="110";
	end if;
	if (ll=239 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=239 and cc>=201 and cc<207) then grbp<="110";
	end if;
	if (ll=239 and cc>=210 and cc<212) then grbp<="110";
	end if;
	if (ll=239 and cc>=213 and cc<216) then grbp<="110";
	end if;
	if (ll=239 and cc>=217 and cc<221) then grbp<="110";
	end if;
	if (cc=245 and ll=239) then grbp<="110";
	end if;
	if (ll=239 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (ll=240 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=138 and ll=240) then grbp<="110";
	end if;
	if (cc=201 and ll=240) then grbp<="110";
	end if;
	if (ll=240 and cc>=201 and cc<216) then grbp<="110";
	end if;
	if (ll=240 and cc>=217 and cc<219) then grbp<="110";
	end if;
	if (cc=242 and ll=240) then grbp<="110";
	end if;
	if (cc=246 and ll=240) then grbp<="110";
	end if;
	if (cc=17 and ll=241) then grbp<="110";
	end if;
	if (ll=241 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=241 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=241 and cc>=199 and cc<208) then grbp<="110";
	end if;
	if (ll=241 and cc>=210 and cc<219) then grbp<="110";
	end if;
	if (cc=242 and ll=241) then grbp<="110";
	end if;
	if (cc=17 and ll=242) then grbp<="110";
	end if;
	if (ll=242 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=199 and ll=242) then grbp<="110";
	end if;
	if (ll=242 and cc>=199 and cc<213) then grbp<="110";
	end if;
	if (ll=242 and cc>=214 and cc<217) then grbp<="110";
	end if;
	if (ll=242 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (cc=232 and ll=242) then grbp<="110";
	end if;
	if (cc=245 and ll=242) then grbp<="110";
	end if;
	if (cc=17 and ll=243) then grbp<="110";
	end if;
	if (ll=243 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=199 and ll=243) then grbp<="110";
	end if;
	if (ll=243 and cc>=199 and cc<210) then grbp<="110";
	end if;
	if (cc=214 and ll=243) then grbp<="110";
	end if;
	if (ll=243 and cc>=214 and cc<217) then grbp<="110";
	end if;
	if (cc=232 and ll=243) then grbp<="110";
	end if;
	if (cc=242 and ll=243) then grbp<="110";
	end if;
	if (cc=17 and ll=244) then grbp<="110";
	end if;
	if (ll=244 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=244 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=199 and ll=244) then grbp<="110";
	end if;
	if (ll=244 and cc>=199 and cc<206) then grbp<="110";
	end if;
	if (ll=244 and cc>=207 and cc<213) then grbp<="110";
	end if;
	if (ll=244 and cc>=214 and cc<218) then grbp<="110";
	end if;
	if (cc=231 and ll=244) then grbp<="110";
	end if;
	if (ll=244 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (cc=242 and ll=244) then grbp<="110";
	end if;
	if (ll=244 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (ll=245 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=245 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (cc=200 and ll=245) then grbp<="110";
	end if;
	if (ll=245 and cc>=200 and cc<210) then grbp<="110";
	end if;
	if (ll=245 and cc>=212 and cc<217) then grbp<="110";
	end if;
	if (cc=220 and ll=245) then grbp<="110";
	end if;
	if (cc=231 and ll=245) then grbp<="110";
	end if;
	if (cc=237 and ll=245) then grbp<="110";
	end if;
	if (ll=245 and cc>=237 and cc<239) then grbp<="110";
	end if;
	if (ll=245 and cc>=242 and cc<244) then grbp<="110";
	end if;
	if (ll=246 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=246 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=138 and ll=246) then grbp<="110";
	end if;
	if (cc=198 and ll=246) then grbp<="110";
	end if;
	if (ll=246 and cc>=198 and cc<205) then grbp<="110";
	end if;
	if (ll=246 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (ll=246 and cc>=209 and cc<212) then grbp<="110";
	end if;
	if (ll=246 and cc>=216 and cc<219) then grbp<="110";
	end if;
	if (cc=238 and ll=246) then grbp<="110";
	end if;
	if (cc=17 and ll=247) then grbp<="110";
	end if;
	if (ll=247 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=137 and ll=247) then grbp<="110";
	end if;
	if (cc=198 and ll=247) then grbp<="110";
	end if;
	if (ll=247 and cc>=198 and cc<209) then grbp<="110";
	end if;
	if (ll=247 and cc>=210 and cc<213) then grbp<="110";
	end if;
	if (cc=218 and ll=247) then grbp<="110";
	end if;
	if (cc=220 and ll=247) then grbp<="110";
	end if;
	if (cc=230 and ll=247) then grbp<="110";
	end if;
	if (cc=234 and ll=247) then grbp<="110";
	end if;
	if (cc=238 and ll=247) then grbp<="110";
	end if;
	if (ll=247 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=248 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (cc=124 and ll=248) then grbp<="110";
	end if;
	if (cc=137 and ll=248) then grbp<="110";
	end if;
	if (cc=198 and ll=248) then grbp<="110";
	end if;
	if (ll=248 and cc>=198 and cc<205) then grbp<="110";
	end if;
	if (ll=248 and cc>=206 and cc<209) then grbp<="110";
	end if;
	if (cc=212 and ll=248) then grbp<="110";
	end if;
	if (ll=248 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=218 and ll=248) then grbp<="110";
	end if;
	if (cc=230 and ll=248) then grbp<="110";
	end if;
	if (cc=238 and ll=248) then grbp<="110";
	end if;
	if (cc=17 and ll=249) then grbp<="110";
	end if;
	if (ll=249 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=249 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (cc=123 and ll=249) then grbp<="110";
	end if;
	if (ll=249 and cc>=123 and cc<125) then grbp<="110";
	end if;
	if (cc=160 and ll=249) then grbp<="110";
	end if;
	if (cc=183 and ll=249) then grbp<="110";
	end if;
	if (cc=197 and ll=249) then grbp<="110";
	end if;
	if (ll=249 and cc>=197 and cc<199) then grbp<="110";
	end if;
	if (ll=249 and cc>=200 and cc<213) then grbp<="110";
	end if;
	if (cc=219 and ll=249) then grbp<="110";
	end if;
	if (cc=229 and ll=249) then grbp<="110";
	end if;
	if (cc=231 and ll=249) then grbp<="110";
	end if;
	if (cc=236 and ll=249) then grbp<="110";
	end if;
	if (ll=249 and cc>=236 and cc<239) then grbp<="110";
	end if;
	if (ll=250 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=124 and ll=250) then grbp<="110";
	end if;
	if (cc=136 and ll=250) then grbp<="110";
	end if;
	if (ll=250 and cc>=136 and cc<139) then grbp<="110";
	end if;
	if (ll=250 and cc>=199 and cc<211) then grbp<="110";
	end if;
	if (cc=229 and ll=250) then grbp<="110";
	end if;
	if (cc=236 and ll=250) then grbp<="110";
	end if;
	if (ll=250 and cc>=236 and cc<238) then grbp<="110";
	end if;
	if (cc=17 and ll=251) then grbp<="110";
	end if;
	if (ll=251 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=136 and ll=251) then grbp<="110";
	end if;
	if (ll=251 and cc>=136 and cc<138) then grbp<="110";
	end if;
	if (cc=200 and ll=251) then grbp<="110";
	end if;
	if (ll=251 and cc>=200 and cc<209) then grbp<="110";
	end if;
	if (cc=215 and ll=251) then grbp<="110";
	end if;
	if (cc=229 and ll=251) then grbp<="110";
	end if;
	if (cc=236 and ll=251) then grbp<="110";
	end if;
	if (cc=238 and ll=251) then grbp<="110";
	end if;
	if (cc=17 and ll=252) then grbp<="110";
	end if;
	if (ll=252 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (ll=252 and cc>=136 and cc<138) then grbp<="110";
	end if;
	if (ll=252 and cc>=197 and cc<209) then grbp<="110";
	end if;
	if (ll=252 and cc>=210 and cc<212) then grbp<="110";
	end if;
	if (cc=228 and ll=252) then grbp<="110";
	end if;
	if (ll=252 and cc>=228 and cc<231) then grbp<="110";
	end if;
	if (cc=235 and ll=252) then grbp<="110";
	end if;
	if (ll=252 and cc>=235 and cc<239) then grbp<="110";
	end if;
	if (ll=253 and cc>=17 and cc<28) then grbp<="110";
	end if;
	if (cc=158 and ll=253) then grbp<="110";
	end if;
	if (cc=197 and ll=253) then grbp<="110";
	end if;
	if (ll=253 and cc>=197 and cc<210) then grbp<="110";
	end if;
	if (ll=253 and cc>=228 and cc<230) then grbp<="110";
	end if;
	if (ll=253 and cc>=233 and cc<236) then grbp<="110";
	end if;
	if (ll=253 and cc>=237 and cc<239) then grbp<="110";
	end if;
	if (ll=254 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=254 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=88 and ll=254) then grbp<="110";
	end if;
	if (cc=101 and ll=254) then grbp<="110";
	end if;
	if (cc=135 and ll=254) then grbp<="110";
	end if;
	if (cc=137 and ll=254) then grbp<="110";
	end if;
	if (cc=159 and ll=254) then grbp<="110";
	end if;
	if (cc=197 and ll=254) then grbp<="110";
	end if;
	if (ll=254 and cc>=197 and cc<212) then grbp<="110";
	end if;
	if (cc=228 and ll=254) then grbp<="110";
	end if;
	if (ll=254 and cc>=228 and cc<230) then grbp<="110";
	end if;
	if (ll=254 and cc>=232 and cc<239) then grbp<="110";
	end if;
	if (ll=255 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=255 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=197 and ll=255) then grbp<="110";
	end if;
	if (ll=255 and cc>=197 and cc<212) then grbp<="110";
	end if;
	if (ll=255 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=255 and cc>=227 and cc<230) then grbp<="110";
	end if;
	if (cc=234 and ll=255) then grbp<="110";
	end if;
	if (ll=255 and cc>=234 and cc<237) then grbp<="110";
	end if;
	if (ll=256 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=256 and cc>=124 and cc<128) then grbp<="110";
	end if;
	if (ll=256 and cc>=135 and cc<137) then grbp<="110";
	end if;
	if (cc=196 and ll=256) then grbp<="110";
	end if;
	if (ll=256 and cc>=196 and cc<210) then grbp<="110";
	end if;
	if (cc=214 and ll=256) then grbp<="110";
	end if;
	if (ll=256 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=256 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=256 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (cc=17 and ll=257) then grbp<="110";
	end if;
	if (ll=257 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=257 and cc>=125 and cc<130) then grbp<="110";
	end if;
	if (cc=135 and ll=257) then grbp<="110";
	end if;
	if (ll=257 and cc>=135 and cc<137) then grbp<="110";
	end if;
	if (cc=196 and ll=257) then grbp<="110";
	end if;
	if (ll=257 and cc>=196 and cc<202) then grbp<="110";
	end if;
	if (ll=257 and cc>=203 and cc<211) then grbp<="110";
	end if;
	if (ll=257 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=257 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=257 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (ll=258 and cc>=17 and cc<19) then grbp<="110";
	end if;
	if (cc=22 and ll=258) then grbp<="110";
	end if;
	if (ll=258 and cc>=22 and cc<29) then grbp<="110";
	end if;
	if (cc=129 and ll=258) then grbp<="110";
	end if;
	if (ll=258 and cc>=129 and cc<132) then grbp<="110";
	end if;
	if (ll=258 and cc>=134 and cc<137) then grbp<="110";
	end if;
	if (ll=258 and cc>=196 and cc<202) then grbp<="110";
	end if;
	if (ll=258 and cc>=203 and cc<212) then grbp<="110";
	end if;
	if (cc=218 and ll=258) then grbp<="110";
	end if;
	if (cc=227 and ll=258) then grbp<="110";
	end if;
	if (ll=258 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=258 and cc>=232 and cc<235) then grbp<="110";
	end if;
	if (ll=259 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=132 and ll=259) then grbp<="110";
	end if;
	if (ll=259 and cc>=132 and cc<137) then grbp<="110";
	end if;
	if (cc=196 and ll=259) then grbp<="110";
	end if;
	if (ll=259 and cc>=196 and cc<215) then grbp<="110";
	end if;
	if (cc=228 and ll=259) then grbp<="110";
	end if;
	if (cc=230 and ll=259) then grbp<="110";
	end if;
	if (ll=259 and cc>=230 and cc<234) then grbp<="110";
	end if;
	if (cc=17 and ll=260) then grbp<="110";
	end if;
	if (ll=260 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=260 and cc>=129 and cc<131) then grbp<="110";
	end if;
	if (cc=135 and ll=260) then grbp<="110";
	end if;
	if (cc=157 and ll=260) then grbp<="110";
	end if;
	if (cc=197 and ll=260) then grbp<="110";
	end if;
	if (ll=260 and cc>=197 and cc<209) then grbp<="110";
	end if;
	if (ll=260 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=226 and ll=260) then grbp<="110";
	end if;
	if (cc=231 and ll=260) then grbp<="110";
	end if;
	if (cc=233 and ll=260) then grbp<="110";
	end if;
	if (cc=17 and ll=261) then grbp<="110";
	end if;
	if (ll=261 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=129 and ll=261) then grbp<="110";
	end if;
	if (cc=135 and ll=261) then grbp<="110";
	end if;
	if (cc=157 and ll=261) then grbp<="110";
	end if;
	if (cc=196 and ll=261) then grbp<="110";
	end if;
	if (ll=261 and cc>=196 and cc<206) then grbp<="110";
	end if;
	if (ll=261 and cc>=207 and cc<211) then grbp<="110";
	end if;
	if (ll=261 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (ll=261 and cc>=215 and cc<217) then grbp<="110";
	end if;
	if (ll=261 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=261 and cc>=231 and cc<233) then grbp<="110";
	end if;
	if (ll=262 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=262 and cc>=79 and cc<81) then grbp<="110";
	end if;
	if (cc=131 and ll=262) then grbp<="110";
	end if;
	if (ll=262 and cc>=131 and cc<133) then grbp<="110";
	end if;
	if (cc=157 and ll=262) then grbp<="110";
	end if;
	if (cc=196 and ll=262) then grbp<="110";
	end if;
	if (ll=262 and cc>=196 and cc<206) then grbp<="110";
	end if;
	if (ll=262 and cc>=207 and cc<213) then grbp<="110";
	end if;
	if (ll=262 and cc>=214 and cc<217) then grbp<="110";
	end if;
	if (ll=262 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=262 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (cc=17 and ll=263) then grbp<="110";
	end if;
	if (ll=263 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=263 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=81 and ll=263) then grbp<="110";
	end if;
	if (cc=131 and ll=263) then grbp<="110";
	end if;
	if (cc=133 and ll=263) then grbp<="110";
	end if;
	if (ll=263 and cc>=133 and cc<135) then grbp<="110";
	end if;
	if (cc=184 and ll=263) then grbp<="110";
	end if;
	if (cc=196 and ll=263) then grbp<="110";
	end if;
	if (ll=263 and cc>=196 and cc<204) then grbp<="110";
	end if;
	if (ll=263 and cc>=205 and cc<211) then grbp<="110";
	end if;
	if (cc=214 and ll=263) then grbp<="110";
	end if;
	if (ll=263 and cc>=214 and cc<218) then grbp<="110";
	end if;
	if (ll=263 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=263 and cc>=229 and cc<234) then grbp<="110";
	end if;
	if (ll=264 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=264 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=127 and ll=264) then grbp<="110";
	end if;
	if (cc=130 and ll=264) then grbp<="110";
	end if;
	if (ll=264 and cc>=130 and cc<134) then grbp<="110";
	end if;
	if (cc=157 and ll=264) then grbp<="110";
	end if;
	if (cc=195 and ll=264) then grbp<="110";
	end if;
	if (ll=264 and cc>=195 and cc<197) then grbp<="110";
	end if;
	if (cc=201 and ll=264) then grbp<="110";
	end if;
	if (ll=264 and cc>=201 and cc<209) then grbp<="110";
	end if;
	if (cc=214 and ll=264) then grbp<="110";
	end if;
	if (ll=264 and cc>=214 and cc<216) then grbp<="110";
	end if;
	if (ll=264 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=264 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (ll=264 and cc>=232 and cc<234) then grbp<="110";
	end if;
	if (ll=265 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=133 and ll=265) then grbp<="110";
	end if;
	if (cc=152 and ll=265) then grbp<="110";
	end if;
	if (cc=195 and ll=265) then grbp<="110";
	end if;
	if (ll=265 and cc>=195 and cc<211) then grbp<="110";
	end if;
	if (ll=265 and cc>=213 and cc<216) then grbp<="110";
	end if;
	if (cc=230 and ll=265) then grbp<="110";
	end if;
	if (cc=232 and ll=265) then grbp<="110";
	end if;
	if (cc=18 and ll=266) then grbp<="110";
	end if;
	if (ll=266 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=266 and cc>=132 and cc<135) then grbp<="110";
	end if;
	if (ll=266 and cc>=196 and cc<203) then grbp<="110";
	end if;
	if (ll=266 and cc>=204 and cc<211) then grbp<="110";
	end if;
	if (ll=266 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (cc=224 and ll=266) then grbp<="110";
	end if;
	if (cc=228 and ll=266) then grbp<="110";
	end if;
	if (cc=230 and ll=266) then grbp<="110";
	end if;
	if (ll=266 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=267 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (ll=267 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=132 and ll=267) then grbp<="110";
	end if;
	if (ll=267 and cc>=132 and cc<135) then grbp<="110";
	end if;
	if (ll=267 and cc>=195 and cc<202) then grbp<="110";
	end if;
	if (ll=267 and cc>=204 and cc<210) then grbp<="110";
	end if;
	if (ll=267 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (cc=230 and ll=267) then grbp<="110";
	end if;
	if (ll=267 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=268 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (ll=268 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (ll=268 and cc>=132 and cc<136) then grbp<="110";
	end if;
	if (cc=196 and ll=268) then grbp<="110";
	end if;
	if (ll=268 and cc>=196 and cc<205) then grbp<="110";
	end if;
	if (ll=268 and cc>=207 and cc<210) then grbp<="110";
	end if;
	if (cc=214 and ll=268) then grbp<="110";
	end if;
	if (cc=216 and ll=268) then grbp<="110";
	end if;
	if (cc=224 and ll=268) then grbp<="110";
	end if;
	if (cc=226 and ll=268) then grbp<="110";
	end if;
	if (ll=268 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (ll=268 and cc>=229 and cc<232) then grbp<="110";
	end if;
	if (ll=269 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=269 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=135 and ll=269) then grbp<="110";
	end if;
	if (cc=195 and ll=269) then grbp<="110";
	end if;
	if (ll=269 and cc>=195 and cc<206) then grbp<="110";
	end if;
	if (ll=269 and cc>=207 and cc<213) then grbp<="110";
	end if;
	if (ll=269 and cc>=224 and cc<227) then grbp<="110";
	end if;
	if (cc=17 and ll=270) then grbp<="110";
	end if;
	if (ll=270 and cc>=17 and cc<20) then grbp<="110";
	end if;
	if (ll=270 and cc>=21 and cc<29) then grbp<="110";
	end if;
	if (ll=270 and cc>=132 and cc<136) then grbp<="110";
	end if;
	if (cc=195 and ll=270) then grbp<="110";
	end if;
	if (ll=270 and cc>=195 and cc<208) then grbp<="110";
	end if;
	if (cc=224 and ll=270) then grbp<="110";
	end if;
	if (ll=270 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (cc=17 and ll=271) then grbp<="110";
	end if;
	if (ll=271 and cc>=17 and cc<20) then grbp<="110";
	end if;
	if (ll=271 and cc>=22 and cc<29) then grbp<="110";
	end if;
	if (ll=271 and cc>=90 and cc<92) then grbp<="110";
	end if;
	if (cc=133 and ll=271) then grbp<="110";
	end if;
	if (ll=271 and cc>=133 and cc<136) then grbp<="110";
	end if;
	if (cc=194 and ll=271) then grbp<="110";
	end if;
	if (ll=271 and cc>=194 and cc<208) then grbp<="110";
	end if;
	if (ll=271 and cc>=209 and cc<211) then grbp<="110";
	end if;
	if (cc=223 and ll=271) then grbp<="110";
	end if;
	if (ll=271 and cc>=223 and cc<226) then grbp<="110";
	end if;
	if (cc=17 and ll=272) then grbp<="110";
	end if;
	if (ll=272 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=272 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=133 and ll=272) then grbp<="110";
	end if;
	if (cc=136 and ll=272) then grbp<="110";
	end if;
	if (cc=194 and ll=272) then grbp<="110";
	end if;
	if (ll=272 and cc>=194 and cc<205) then grbp<="110";
	end if;
	if (ll=272 and cc>=206 and cc<210) then grbp<="110";
	end if;
	if (cc=213 and ll=272) then grbp<="110";
	end if;
	if (cc=223 and ll=272) then grbp<="110";
	end if;
	if (ll=272 and cc>=223 and cc<226) then grbp<="110";
	end if;
	if (ll=272 and cc>=227 and cc<230) then grbp<="110";
	end if;
	if (ll=273 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=273 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=135 and ll=273) then grbp<="110";
	end if;
	if (ll=273 and cc>=135 and cc<138) then grbp<="110";
	end if;
	if (ll=273 and cc>=194 and cc<207) then grbp<="110";
	end if;
	if (cc=223 and ll=273) then grbp<="110";
	end if;
	if (ll=273 and cc>=223 and cc<225) then grbp<="110";
	end if;
	if (cc=228 and ll=273) then grbp<="110";
	end if;
	if (cc=16 and ll=274) then grbp<="110";
	end if;
	if (ll=274 and cc>=16 and cc<29) then grbp<="110";
	end if;
	if (cc=93 and ll=274) then grbp<="110";
	end if;
	if (cc=134 and ll=274) then grbp<="110";
	end if;
	if (cc=194 and ll=274) then grbp<="110";
	end if;
	if (ll=274 and cc>=194 and cc<206) then grbp<="110";
	end if;
	if (ll=274 and cc>=207 and cc<210) then grbp<="110";
	end if;
	if (ll=274 and cc>=223 and cc<226) then grbp<="110";
	end if;
	if (cc=17 and ll=275) then grbp<="110";
	end if;
	if (ll=275 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=275 and cc>=133 and cc<135) then grbp<="110";
	end if;
	if (cc=147 and ll=275) then grbp<="110";
	end if;
	if (cc=194 and ll=275) then grbp<="110";
	end if;
	if (ll=275 and cc>=194 and cc<203) then grbp<="110";
	end if;
	if (ll=275 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (ll=275 and cc>=208 and cc<211) then grbp<="110";
	end if;
	if (ll=275 and cc>=223 and cc<226) then grbp<="110";
	end if;
	if (cc=16 and ll=276) then grbp<="110";
	end if;
	if (ll=276 and cc>=16 and cc<29) then grbp<="110";
	end if;
	if (ll=276 and cc>=133 and cc<135) then grbp<="110";
	end if;
	if (cc=193 and ll=276) then grbp<="110";
	end if;
	if (ll=276 and cc>=193 and cc<205) then grbp<="110";
	end if;
	if (cc=210 and ll=276) then grbp<="110";
	end if;
	if (cc=214 and ll=276) then grbp<="110";
	end if;
	if (cc=223 and ll=276) then grbp<="110";
	end if;
	if (ll=276 and cc>=223 and cc<229) then grbp<="110";
	end if;
	if (ll=277 and cc>=16 and cc<23) then grbp<="110";
	end if;
	if (ll=277 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=156 and ll=277) then grbp<="110";
	end if;
	if (cc=194 and ll=277) then grbp<="110";
	end if;
	if (ll=277 and cc>=194 and cc<207) then grbp<="110";
	end if;
	if (cc=213 and ll=277) then grbp<="110";
	end if;
	if (ll=277 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (ll=277 and cc>=223 and cc<225) then grbp<="110";
	end if;
	if (ll=277 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (ll=278 and cc>=16 and cc<25) then grbp<="110";
	end if;
	if (ll=278 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=190 and ll=278) then grbp<="110";
	end if;
	if (cc=193 and ll=278) then grbp<="110";
	end if;
	if (ll=278 and cc>=193 and cc<206) then grbp<="110";
	end if;
	if (ll=278 and cc>=207 and cc<209) then grbp<="110";
	end if;
	if (ll=278 and cc>=223 and cc<228) then grbp<="110";
	end if;
	if (ll=279 and cc>=16 and cc<29) then grbp<="110";
	end if;
	if (cc=193 and ll=279) then grbp<="110";
	end if;
	if (ll=279 and cc>=193 and cc<203) then grbp<="110";
	end if;
	if (cc=206 and ll=279) then grbp<="110";
	end if;
	if (cc=209 and ll=279) then grbp<="110";
	end if;
	if (cc=215 and ll=279) then grbp<="110";
	end if;
	if (cc=223 and ll=279) then grbp<="110";
	end if;
	if (ll=279 and cc>=223 and cc<228) then grbp<="110";
	end if;
	if (ll=280 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=280 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=136 and ll=280) then grbp<="110";
	end if;
	if (cc=156 and ll=280) then grbp<="110";
	end if;
	if (cc=193 and ll=280) then grbp<="110";
	end if;
	if (ll=280 and cc>=193 and cc<205) then grbp<="110";
	end if;
	if (ll=280 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (cc=222 and ll=280) then grbp<="110";
	end if;
	if (ll=280 and cc>=222 and cc<227) then grbp<="110";
	end if;
	if (ll=281 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=281 and cc>=193 and cc<203) then grbp<="110";
	end if;
	if (cc=206 and ll=281) then grbp<="110";
	end if;
	if (ll=281 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (ll=281 and cc>=222 and cc<227) then grbp<="110";
	end if;
	if (ll=282 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=282 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (ll=282 and cc>=193 and cc<201) then grbp<="110";
	end if;
	if (cc=205 and ll=282) then grbp<="110";
	end if;
	if (ll=282 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (cc=213 and ll=282) then grbp<="110";
	end if;
	if (cc=222 and ll=282) then grbp<="110";
	end if;
	if (ll=282 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (cc=16 and ll=283) then grbp<="110";
	end if;
	if (ll=283 and cc>=16 and cc<29) then grbp<="110";
	end if;
	if (cc=193 and ll=283) then grbp<="110";
	end if;
	if (ll=283 and cc>=193 and cc<205) then grbp<="110";
	end if;
	if (cc=209 and ll=283) then grbp<="110";
	end if;
	if (cc=213 and ll=283) then grbp<="110";
	end if;
	if (cc=222 and ll=283) then grbp<="110";
	end if;
	if (ll=283 and cc>=222 and cc<227) then grbp<="110";
	end if;
	if (ll=284 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (ll=284 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=284 and cc>=192 and cc<203) then grbp<="110";
	end if;
	if (cc=209 and ll=284) then grbp<="110";
	end if;
	if (cc=212 and ll=284) then grbp<="110";
	end if;
	if (cc=222 and ll=284) then grbp<="110";
	end if;
	if (ll=284 and cc>=222 and cc<226) then grbp<="110";
	end if;
	if (ll=285 and cc>=16 and cc<24) then grbp<="110";
	end if;
	if (ll=285 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=192 and ll=285) then grbp<="110";
	end if;
	if (ll=285 and cc>=192 and cc<202) then grbp<="110";
	end if;
	if (cc=206 and ll=285) then grbp<="110";
	end if;
	if (cc=209 and ll=285) then grbp<="110";
	end if;
	if (cc=222 and ll=285) then grbp<="110";
	end if;
	if (ll=285 and cc>=222 and cc<225) then grbp<="110";
	end if;
	if (ll=286 and cc>=16 and cc<24) then grbp<="110";
	end if;
	if (ll=286 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (ll=286 and cc>=142 and cc<146) then grbp<="110";
	end if;
	if (cc=192 and ll=286) then grbp<="110";
	end if;
	if (ll=286 and cc>=192 and cc<202) then grbp<="110";
	end if;
	if (ll=286 and cc>=203 and cc<208) then grbp<="110";
	end if;
	if (ll=286 and cc>=222 and cc<226) then grbp<="110";
	end if;
	if (ll=287 and cc>=16 and cc<25) then grbp<="110";
	end if;
	if (ll=287 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=149 and ll=287) then grbp<="110";
	end if;
	if (cc=192 and ll=287) then grbp<="110";
	end if;
	if (ll=287 and cc>=192 and cc<201) then grbp<="110";
	end if;
	if (ll=287 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (ll=287 and cc>=208 and cc<210) then grbp<="110";
	end if;
	if (ll=287 and cc>=222 and cc<225) then grbp<="110";
	end if;
	if (ll=288 and cc>=16 and cc<22) then grbp<="110";
	end if;
	if (ll=288 and cc>=23 and cc<26) then grbp<="110";
	end if;
	if (ll=288 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=192 and ll=288) then grbp<="110";
	end if;
	if (ll=288 and cc>=192 and cc<201) then grbp<="110";
	end if;
	if (ll=288 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (ll=288 and cc>=207 and cc<209) then grbp<="110";
	end if;
	if (cc=222 and ll=288) then grbp<="110";
	end if;
	if (ll=288 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (cc=18 and ll=289) then grbp<="110";
	end if;
	if (ll=289 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (cc=25 and ll=289) then grbp<="110";
	end if;
	if (ll=289 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=192 and ll=289) then grbp<="110";
	end if;
	if (ll=289 and cc>=192 and cc<203) then grbp<="110";
	end if;
	if (ll=289 and cc>=204 and cc<207) then grbp<="110";
	end if;
	if (cc=222 and ll=289) then grbp<="110";
	end if;
	if (ll=289 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=290 and cc>=16 and cc<23) then grbp<="110";
	end if;
	if (ll=290 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=290 and cc>=192 and cc<203) then grbp<="110";
	end if;
	if (ll=290 and cc>=204 and cc<207) then grbp<="110";
	end if;
	if (ll=290 and cc>=209 and cc<211) then grbp<="110";
	end if;
	if (ll=290 and cc>=222 and cc<225) then grbp<="110";
	end if;
	if (ll=291 and cc>=17 and cc<23) then grbp<="110";
	end if;
	if (ll=291 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=291 and cc>=192 and cc<194) then grbp<="110";
	end if;
	if (ll=291 and cc>=195 and cc<202) then grbp<="110";
	end if;
	if (ll=291 and cc>=203 and cc<207) then grbp<="110";
	end if;
	if (ll=291 and cc>=208 and cc<210) then grbp<="110";
	end if;
	if (ll=291 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=292 and cc>=16 and cc<19) then grbp<="110";
	end if;
	if (cc=22 and ll=292) then grbp<="110";
	end if;
	if (ll=292 and cc>=22 and cc<29) then grbp<="110";
	end if;
	if (cc=188 and ll=292) then grbp<="110";
	end if;
	if (cc=192 and ll=292) then grbp<="110";
	end if;
	if (ll=292 and cc>=192 and cc<203) then grbp<="110";
	end if;
	if (ll=292 and cc>=204 and cc<206) then grbp<="110";
	end if;
	if (ll=292 and cc>=207 and cc<210) then grbp<="110";
	end if;
	if (cc=16 and ll=293) then grbp<="110";
	end if;
	if (ll=293 and cc>=16 and cc<21) then grbp<="110";
	end if;
	if (ll=293 and cc>=22 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=293) then grbp<="110";
	end if;
	if (ll=293 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=191 and ll=293) then grbp<="110";
	end if;
	if (ll=293 and cc>=191 and cc<204) then grbp<="110";
	end if;
	if (ll=293 and cc>=207 and cc<209) then grbp<="110";
	end if;
	if (cc=17 and ll=294) then grbp<="110";
	end if;
	if (ll=294 and cc>=17 and cc<21) then grbp<="110";
	end if;
	if (ll=294 and cc>=22 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=294) then grbp<="110";
	end if;
	if (ll=294 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=191 and ll=294) then grbp<="110";
	end if;
	if (ll=294 and cc>=191 and cc<203) then grbp<="110";
	end if;
	if (cc=208 and ll=294) then grbp<="110";
	end if;
	if (cc=210 and ll=294) then grbp<="110";
	end if;
	if (cc=222 and ll=294) then grbp<="110";
	end if;
	if (cc=16 and ll=295) then grbp<="110";
	end if;
	if (ll=295 and cc>=16 and cc<24) then grbp<="110";
	end if;
	if (ll=295 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (ll=295 and cc>=191 and cc<209) then grbp<="110";
	end if;
	if (cc=222 and ll=295) then grbp<="110";
	end if;
	if (cc=16 and ll=296) then grbp<="110";
	end if;
	if (ll=296 and cc>=16 and cc<21) then grbp<="110";
	end if;
	if (cc=24 and ll=296) then grbp<="110";
	end if;
	if (ll=296 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (cc=188 and ll=296) then grbp<="110";
	end if;
	if (cc=190 and ll=296) then grbp<="110";
	end if;
	if (ll=296 and cc>=190 and cc<207) then grbp<="110";
	end if;
	if (cc=212 and ll=296) then grbp<="110";
	end if;
	if (cc=222 and ll=296) then grbp<="110";
	end if;
	if (cc=17 and ll=297) then grbp<="110";
	end if;
	if (ll=297 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=297 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=297 and cc>=81 and cc<83) then grbp<="110";
	end if;
	if (cc=190 and ll=297) then grbp<="110";
	end if;
	if (ll=297 and cc>=190 and cc<209) then grbp<="110";
	end if;
	if (cc=222 and ll=297) then grbp<="110";
	end if;
	if (cc=17 and ll=298) then grbp<="110";
	end if;
	if (ll=298 and cc>=17 and cc<21) then grbp<="110";
	end if;
	if (ll=298 and cc>=22 and cc<27) then grbp<="110";
	end if;
	if (cc=187 and ll=298) then grbp<="110";
	end if;
	if (ll=298 and cc>=187 and cc<189) then grbp<="110";
	end if;
	if (ll=298 and cc>=192 and cc<209) then grbp<="110";
	end if;
	if (cc=16 and ll=299) then grbp<="110";
	end if;
	if (ll=299 and cc>=16 and cc<25) then grbp<="110";
	end if;
	if (cc=188 and ll=299) then grbp<="110";
	end if;
	if (cc=190 and ll=299) then grbp<="110";
	end if;
	if (ll=299 and cc>=190 and cc<208) then grbp<="110";
	end if;
	if (ll=299 and cc>=211 and cc<213) then grbp<="110";
	end if;
	if (cc=16 and ll=300) then grbp<="110";
	end if;
	if (ll=300 and cc>=16 and cc<26) then grbp<="110";
	end if;
	if (cc=80 and ll=300) then grbp<="110";
	end if;
	if (cc=188 and ll=300) then grbp<="110";
	end if;
	if (cc=190 and ll=300) then grbp<="110";
	end if;
	if (ll=300 and cc>=190 and cc<209) then grbp<="110";
	end if;
	if (cc=17 and ll=301) then grbp<="110";
	end if;
	if (ll=301 and cc>=17 and cc<20) then grbp<="110";
	end if;
	if (cc=23 and ll=301) then grbp<="110";
	end if;
	if (ll=301 and cc>=23 and cc<26) then grbp<="110";
	end if;
	if (ll=301 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=81 and ll=301) then grbp<="110";
	end if;
	if (cc=188 and ll=301) then grbp<="110";
	end if;
	if (cc=190 and ll=301) then grbp<="110";
	end if;
	if (ll=301 and cc>=190 and cc<209) then grbp<="110";
	end if;
	if (ll=302 and cc>=17 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=302) then grbp<="110";
	end if;
	if (ll=302 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (ll=302 and cc>=78 and cc<80) then grbp<="110";
	end if;
	if (cc=190 and ll=302) then grbp<="110";
	end if;
	if (ll=302 and cc>=190 and cc<210) then grbp<="110";
	end if;
	if (cc=222 and ll=302) then grbp<="110";
	end if;
	if (cc=17 and ll=303) then grbp<="110";
	end if;
	if (ll=303 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=303 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (ll=303 and cc>=78 and cc<80) then grbp<="110";
	end if;
	if (cc=191 and ll=303) then grbp<="110";
	end if;
	if (ll=303 and cc>=191 and cc<209) then grbp<="110";
	end if;
	if (ll=304 and cc>=17 and cc<26) then grbp<="110";
	end if;
	if (ll=304 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=188 and ll=304) then grbp<="110";
	end if;
	if (cc=190 and ll=304) then grbp<="110";
	end if;
	if (ll=304 and cc>=190 and cc<207) then grbp<="110";
	end if;
	if (ll=304 and cc>=208 and cc<210) then grbp<="110";
	end if;
	if (ll=305 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=186 and ll=305) then grbp<="110";
	end if;
	if (cc=188 and ll=305) then grbp<="110";
	end if;
	if (cc=190 and ll=305) then grbp<="110";
	end if;
	if (ll=305 and cc>=190 and cc<212) then grbp<="110";
	end if;
	if (ll=306 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=187 and ll=306) then grbp<="110";
	end if;
	if (cc=190 and ll=306) then grbp<="110";
	end if;
	if (ll=306 and cc>=190 and cc<200) then grbp<="110";
	end if;
	if (ll=306 and cc>=201 and cc<211) then grbp<="110";
	end if;
	if (cc=20 and ll=307) then grbp<="110";
	end if;
	if (ll=307 and cc>=20 and cc<25) then grbp<="110";
	end if;
	if (ll=307 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (ll=307 and cc>=144 and cc<146) then grbp<="110";
	end if;
	if (cc=190 and ll=307) then grbp<="110";
	end if;
	if (ll=307 and cc>=190 and cc<197) then grbp<="110";
	end if;
	if (ll=307 and cc>=198 and cc<210) then grbp<="110";
	end if;
	if (ll=307 and cc>=211 and cc<213) then grbp<="110";
	end if;
	if (ll=308 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=308 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=145 and ll=308) then grbp<="110";
	end if;
	if (ll=308 and cc>=145 and cc<147) then grbp<="110";
	end if;
	if (cc=190 and ll=308) then grbp<="110";
	end if;
	if (ll=308 and cc>=190 and cc<198) then grbp<="110";
	end if;
	if (ll=308 and cc>=199 and cc<204) then grbp<="110";
	end if;
	if (ll=308 and cc>=205 and cc<209) then grbp<="110";
	end if;
	if (cc=18 and ll=309) then grbp<="110";
	end if;
	if (ll=309 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=189 and ll=309) then grbp<="110";
	end if;
	if (ll=309 and cc>=189 and cc<199) then grbp<="110";
	end if;
	if (ll=309 and cc>=200 and cc<204) then grbp<="110";
	end if;
	if (ll=309 and cc>=205 and cc<210) then grbp<="110";
	end if;
	if (cc=18 and ll=310) then grbp<="110";
	end if;
	if (ll=310 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=310 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=189 and ll=310) then grbp<="110";
	end if;
	if (ll=310 and cc>=189 and cc<195) then grbp<="110";
	end if;
	if (cc=198 and ll=310) then grbp<="110";
	end if;
	if (ll=310 and cc>=198 and cc<210) then grbp<="110";
	end if;
	if (cc=221 and ll=310) then grbp<="110";
	end if;
	if (cc=18 and ll=311) then grbp<="110";
	end if;
	if (ll=311 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=190 and ll=311) then grbp<="110";
	end if;
	if (ll=311 and cc>=190 and cc<211) then grbp<="110";
	end if;
	if (cc=18 and ll=312) then grbp<="110";
	end if;
	if (ll=312 and cc>=18 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=312) then grbp<="110";
	end if;
	if (ll=312 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=190 and ll=312) then grbp<="110";
	end if;
	if (ll=312 and cc>=190 and cc<195) then grbp<="110";
	end if;
	if (ll=312 and cc>=197 and cc<200) then grbp<="110";
	end if;
	if (ll=312 and cc>=201 and cc<209) then grbp<="110";
	end if;
	if (ll=313 and cc>=18 and cc<24) then grbp<="110";
	end if;
	if (ll=313 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (cc=187 and ll=313) then grbp<="110";
	end if;
	if (cc=189 and ll=313) then grbp<="110";
	end if;
	if (ll=313 and cc>=189 and cc<192) then grbp<="110";
	end if;
	if (ll=313 and cc>=193 and cc<200) then grbp<="110";
	end if;
	if (ll=313 and cc>=201 and cc<206) then grbp<="110";
	end if;
	if (cc=209 and ll=313) then grbp<="110";
	end if;
	if (cc=221 and ll=313) then grbp<="110";
	end if;
	if (cc=17 and ll=314) then grbp<="110";
	end if;
	if (ll=314 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=189 and ll=314) then grbp<="110";
	end if;
	if (ll=314 and cc>=189 and cc<192) then grbp<="110";
	end if;
	if (ll=314 and cc>=193 and cc<199) then grbp<="110";
	end if;
	if (ll=314 and cc>=200 and cc<210) then grbp<="110";
	end if;
	if (ll=315 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=315 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (ll=315 and cc>=189 and cc<196) then grbp<="110";
	end if;
	if (ll=315 and cc>=197 and cc<200) then grbp<="110";
	end if;
	if (ll=315 and cc>=201 and cc<208) then grbp<="110";
	end if;
	if (ll=315 and cc>=249 and cc<251) then grbp<="110";
	end if;
	if (ll=316 and cc>=17 and cc<21) then grbp<="110";
	end if;
	if (ll=316 and cc>=22 and cc<29) then grbp<="110";
	end if;
	if (cc=189 and ll=316) then grbp<="110";
	end if;
	if (ll=316 and cc>=189 and cc<197) then grbp<="110";
	end if;
	if (ll=316 and cc>=198 and cc<200) then grbp<="110";
	end if;
	if (ll=316 and cc>=202 and cc<205) then grbp<="110";
	end if;
	if (ll=316 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (cc=247 and ll=316) then grbp<="110";
	end if;
	if (ll=316 and cc>=247 and cc<249) then grbp<="110";
	end if;
	if (ll=317 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=317 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=193 and ll=317) then grbp<="110";
	end if;
	if (ll=317 and cc>=193 and cc<197) then grbp<="110";
	end if;
	if (cc=201 and ll=317) then grbp<="110";
	end if;
	if (ll=317 and cc>=201 and cc<203) then grbp<="110";
	end if;
	if (ll=317 and cc>=205 and cc<207) then grbp<="110";
	end if;
	if (ll=317 and cc>=245 and cc<247) then grbp<="110";
	end if;
	if (ll=318 and cc>=18 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=318) then grbp<="110";
	end if;
	if (ll=318 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=186 and ll=318) then grbp<="110";
	end if;
	if (ll=318 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=200 and ll=318) then grbp<="110";
	end if;
	if (ll=318 and cc>=200 and cc<208) then grbp<="110";
	end if;
	if (cc=244 and ll=318) then grbp<="110";
	end if;
	if (ll=318 and cc>=244 and cc<246) then grbp<="110";
	end if;
	if (ll=319 and cc>=17 and cc<22) then grbp<="110";
	end if;
	if (ll=319 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (ll=319 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=200 and ll=319) then grbp<="110";
	end if;
	if (ll=319 and cc>=200 and cc<202) then grbp<="110";
	end if;
	if (ll=319 and cc>=203 and cc<208) then grbp<="110";
	end if;
	if (cc=242 and ll=319) then grbp<="110";
	end if;
	if (ll=319 and cc>=242 and cc<245) then grbp<="110";
	end if;
	if (ll=320 and cc>=17 and cc<25) then grbp<="110";
	end if;
	if (ll=320 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (cc=200 and ll=320) then grbp<="110";
	end if;
	if (ll=320 and cc>=200 and cc<205) then grbp<="110";
	end if;
	if (cc=220 and ll=320) then grbp<="110";
	end if;
	if (cc=241 and ll=320) then grbp<="110";
	end if;
	if (ll=320 and cc>=241 and cc<243) then grbp<="110";
	end if;
	if (ll=321 and cc>=17 and cc<20) then grbp<="110";
	end if;
	if (ll=321 and cc>=21 and cc<26) then grbp<="110";
	end if;
	if (ll=321 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=204 and ll=321) then grbp<="110";
	end if;
	if (cc=206 and ll=321) then grbp<="110";
	end if;
	if (cc=241 and ll=321) then grbp<="110";
	end if;
	if (cc=17 and ll=322) then grbp<="110";
	end if;
	if (ll=322 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=137 and ll=322) then grbp<="110";
	end if;
	if (cc=139 and ll=322) then grbp<="110";
	end if;
	if (cc=186 and ll=322) then grbp<="110";
	end if;
	if (cc=204 and ll=322) then grbp<="110";
	end if;
	if (ll=322 and cc>=204 and cc<207) then grbp<="110";
	end if;
	if (ll=322 and cc>=239 and cc<241) then grbp<="110";
	end if;
	if (ll=323 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (ll=323 and cc>=137 and cc<139) then grbp<="110";
	end if;
	if (ll=323 and cc>=140 and cc<143) then grbp<="110";
	end if;
	if (cc=239 and ll=323) then grbp<="110";
	end if;
	if (cc=17 and ll=324) then grbp<="110";
	end if;
	if (ll=324 and cc>=17 and cc<19) then grbp<="110";
	end if;
	if (ll=324 and cc>=20 and cc<29) then grbp<="110";
	end if;
	if (cc=142 and ll=324) then grbp<="110";
	end if;
	if (ll=324 and cc>=142 and cc<145) then grbp<="110";
	end if;
	if (cc=184 and ll=324) then grbp<="110";
	end if;
	if (ll=324 and cc>=184 and cc<187) then grbp<="110";
	end if;
	if (ll=324 and cc>=238 and cc<240) then grbp<="110";
	end if;
	if (ll=325 and cc>=17 and cc<29) then grbp<="110";
	end if;
	if (cc=184 and ll=325) then grbp<="110";
	end if;
	if (ll=325 and cc>=184 and cc<187) then grbp<="110";
	end if;
	if (cc=18 and ll=326) then grbp<="110";
	end if;
	if (ll=326 and cc>=18 and cc<23) then grbp<="110";
	end if;
	if (ll=326 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (cc=238 and ll=326) then grbp<="110";
	end if;
	if (cc=18 and ll=327) then grbp<="110";
	end if;
	if (ll=327 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (cc=24 and ll=327) then grbp<="110";
	end if;
	if (ll=327 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (cc=18 and ll=328) then grbp<="110";
	end if;
	if (ll=328 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=237 and ll=328) then grbp<="110";
	end if;
	if (cc=18 and ll=329) then grbp<="110";
	end if;
	if (ll=329 and cc>=18 and cc<28) then grbp<="110";
	end if;
	if (cc=185 and ll=329) then grbp<="110";
	end if;
	if (cc=236 and ll=329) then grbp<="110";
	end if;
	if (cc=18 and ll=330) then grbp<="110";
	end if;
	if (ll=330 and cc>=18 and cc<26) then grbp<="110";
	end if;
	if (cc=235 and ll=330) then grbp<="110";
	end if;
	if (ll=330 and cc>=235 and cc<237) then grbp<="110";
	end if;
	if (ll=331 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (cc=145 and ll=331) then grbp<="110";
	end if;
	if (cc=185 and ll=331) then grbp<="110";
	end if;
	if (cc=220 and ll=331) then grbp<="110";
	end if;
	if (cc=235 and ll=331) then grbp<="110";
	end if;
	if (cc=18 and ll=332) then grbp<="110";
	end if;
	if (cc=20 and ll=332) then grbp<="110";
	end if;
	if (cc=22 and ll=332) then grbp<="110";
	end if;
	if (ll=332 and cc>=22 and cc<25) then grbp<="110";
	end if;
	if (ll=332 and cc>=28 and cc<30) then grbp<="110";
	end if;
	if (cc=220 and ll=332) then grbp<="110";
	end if;
	if (cc=235 and ll=332) then grbp<="110";
	end if;
	if (cc=18 and ll=333) then grbp<="110";
	end if;
	if (ll=333 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=333 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=233 and ll=333) then grbp<="110";
	end if;
	if (ll=333 and cc>=233 and cc<235) then grbp<="110";
	end if;
	if (ll=334 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=189 and ll=334) then grbp<="110";
	end if;
	if (cc=233 and ll=334) then grbp<="110";
	end if;
	if (cc=18 and ll=335) then grbp<="110";
	end if;
	if (ll=335 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=232 and ll=335) then grbp<="110";
	end if;
	if (cc=18 and ll=336) then grbp<="110";
	end if;
	if (ll=336 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=336 and cc>=143 and cc<145) then grbp<="110";
	end if;
	if (cc=191 and ll=336) then grbp<="110";
	end if;
	if (cc=232 and ll=336) then grbp<="110";
	end if;
	if (cc=18 and ll=337) then grbp<="110";
	end if;
	if (ll=337 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=337 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=337 and cc>=143 and cc<145) then grbp<="110";
	end if;
	if (cc=187 and ll=337) then grbp<="110";
	end if;
	if (cc=190 and ll=337) then grbp<="110";
	end if;
	if (cc=231 and ll=337) then grbp<="110";
	end if;
	if (cc=18 and ll=338) then grbp<="110";
	end if;
	if (ll=338 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (ll=338 and cc>=21 and cc<29) then grbp<="110";
	end if;
	if (ll=338 and cc>=142 and cc<144) then grbp<="110";
	end if;
	if (cc=184 and ll=338) then grbp<="110";
	end if;
	if (cc=187 and ll=338) then grbp<="110";
	end if;
	if (cc=190 and ll=338) then grbp<="110";
	end if;
	if (cc=219 and ll=338) then grbp<="110";
	end if;
	if (cc=231 and ll=338) then grbp<="110";
	end if;
	if (cc=18 and ll=339) then grbp<="110";
	end if;
	if (ll=339 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=339 and cc>=142 and cc<145) then grbp<="110";
	end if;
	if (cc=187 and ll=339) then grbp<="110";
	end if;
	if (cc=189 and ll=339) then grbp<="110";
	end if;
	if (cc=219 and ll=339) then grbp<="110";
	end if;
	if (cc=231 and ll=339) then grbp<="110";
	end if;
	if (cc=18 and ll=340) then grbp<="110";
	end if;
	if (ll=340 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=340 and cc>=143 and cc<146) then grbp<="110";
	end if;
	if (cc=187 and ll=340) then grbp<="110";
	end if;
	if (ll=340 and cc>=187 and cc<189) then grbp<="110";
	end if;
	if (cc=219 and ll=340) then grbp<="110";
	end if;
	if (cc=231 and ll=340) then grbp<="110";
	end if;
	if (cc=18 and ll=341) then grbp<="110";
	end if;
	if (ll=341 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (cc=187 and ll=341) then grbp<="110";
	end if;
	if (ll=341 and cc>=187 and cc<189) then grbp<="110";
	end if;
	if (cc=230 and ll=341) then grbp<="110";
	end if;
	if (ll=341 and cc>=230 and cc<232) then grbp<="110";
	end if;
	if (ll=342 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=342 and cc>=142 and cc<145) then grbp<="110";
	end if;
	if (cc=187 and ll=342) then grbp<="110";
	end if;
	if (cc=189 and ll=342) then grbp<="110";
	end if;
	if (ll=342 and cc>=189 and cc<192) then grbp<="110";
	end if;
	if (ll=342 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (ll=343 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=343 and cc>=142 and cc<146) then grbp<="110";
	end if;
	if (cc=187 and ll=343) then grbp<="110";
	end if;
	if (ll=343 and cc>=187 and cc<193) then grbp<="110";
	end if;
	if (ll=343 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (ll=344 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (ll=344 and cc>=22 and cc<29) then grbp<="110";
	end if;
	if (ll=344 and cc>=142 and cc<147) then grbp<="110";
	end if;
	if (ll=344 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (cc=218 and ll=344) then grbp<="110";
	end if;
	if (cc=229 and ll=344) then grbp<="110";
	end if;
	if (ll=344 and cc>=229 and cc<231) then grbp<="110";
	end if;
	if (ll=345 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=345 and cc>=143 and cc<148) then grbp<="110";
	end if;
	if (ll=345 and cc>=187 and cc<192) then grbp<="110";
	end if;
	if (cc=229 and ll=345) then grbp<="110";
	end if;
	if (cc=18 and ll=346) then grbp<="110";
	end if;
	if (ll=346 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (ll=346 and cc>=21 and cc<29) then grbp<="110";
	end if;
	if (ll=346 and cc>=143 and cc<149) then grbp<="110";
	end if;
	if (cc=191 and ll=346) then grbp<="110";
	end if;
	if (cc=218 and ll=346) then grbp<="110";
	end if;
	if (cc=229 and ll=346) then grbp<="110";
	end if;
	if (cc=18 and ll=347) then grbp<="110";
	end if;
	if (ll=347 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (ll=347 and cc>=22 and cc<30) then grbp<="110";
	end if;
	if (ll=347 and cc>=143 and cc<149) then grbp<="110";
	end if;
	if (ll=347 and cc>=189 and cc<191) then grbp<="110";
	end if;
	if (cc=218 and ll=347) then grbp<="110";
	end if;
	if (cc=229 and ll=347) then grbp<="110";
	end if;
	if (cc=18 and ll=348) then grbp<="110";
	end if;
	if (ll=348 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=348 and cc>=144 and cc<149) then grbp<="110";
	end if;
	if (cc=187 and ll=348) then grbp<="110";
	end if;
	if (cc=218 and ll=348) then grbp<="110";
	end if;
	if (cc=18 and ll=349) then grbp<="110";
	end if;
	if (ll=349 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=349 and cc>=143 and cc<149) then grbp<="110";
	end if;
	if (cc=187 and ll=349) then grbp<="110";
	end if;
	if (ll=349 and cc>=187 and cc<189) then grbp<="110";
	end if;
	if (ll=349 and cc>=217 and cc<219) then grbp<="110";
	end if;
	if (cc=18 and ll=350) then grbp<="110";
	end if;
	if (ll=350 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (cc=23 and ll=350) then grbp<="110";
	end if;
	if (cc=25 and ll=350) then grbp<="110";
	end if;
	if (ll=350 and cc>=25 and cc<29) then grbp<="110";
	end if;
	if (ll=350 and cc>=144 and cc<147) then grbp<="110";
	end if;
	if (ll=350 and cc>=148 and cc<150) then grbp<="110";
	end if;
	if (cc=187 and ll=350) then grbp<="110";
	end if;
	if (cc=215 and ll=350) then grbp<="110";
	end if;
	if (ll=350 and cc>=215 and cc<219) then grbp<="110";
	end if;
	if (cc=18 and ll=351) then grbp<="110";
	end if;
	if (ll=351 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=351 and cc>=144 and cc<148) then grbp<="110";
	end if;
	if (cc=183 and ll=351) then grbp<="110";
	end if;
	if (cc=186 and ll=351) then grbp<="110";
	end if;
	if (cc=189 and ll=351) then grbp<="110";
	end if;
	if (cc=214 and ll=351) then grbp<="110";
	end if;
	if (ll=351 and cc>=214 and cc<218) then grbp<="110";
	end if;
	if (cc=18 and ll=352) then grbp<="110";
	end if;
	if (ll=352 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=352 and cc>=145 and cc<149) then grbp<="110";
	end if;
	if (cc=186 and ll=352) then grbp<="110";
	end if;
	if (ll=352 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=214 and ll=352) then grbp<="110";
	end if;
	if (ll=352 and cc>=214 and cc<217) then grbp<="110";
	end if;
	if (ll=352 and cc>=227 and cc<229) then grbp<="110";
	end if;
	if (ll=353 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=353 and cc>=145 and cc<149) then grbp<="110";
	end if;
	if (cc=186 and ll=353) then grbp<="110";
	end if;
	if (ll=353 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=213 and ll=353) then grbp<="110";
	end if;
	if (ll=353 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=18 and ll=354) then grbp<="110";
	end if;
	if (ll=354 and cc>=18 and cc<26) then grbp<="110";
	end if;
	if (ll=354 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (ll=354 and cc>=144 and cc<150) then grbp<="110";
	end if;
	if (ll=354 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (ll=354 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=18 and ll=355) then grbp<="110";
	end if;
	if (ll=355 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (cc=24 and ll=355) then grbp<="110";
	end if;
	if (ll=355 and cc>=24 and cc<30) then grbp<="110";
	end if;
	if (ll=355 and cc>=144 and cc<149) then grbp<="110";
	end if;
	if (cc=183 and ll=355) then grbp<="110";
	end if;
	if (cc=186 and ll=355) then grbp<="110";
	end if;
	if (ll=355 and cc>=186 and cc<190) then grbp<="110";
	end if;
	if (cc=212 and ll=355) then grbp<="110";
	end if;
	if (ll=355 and cc>=212 and cc<214) then grbp<="110";
	end if;
	if (ll=355 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (ll=356 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (ll=356 and cc>=22 and cc<30) then grbp<="110";
	end if;
	if (cc=146 and ll=356) then grbp<="110";
	end if;
	if (ll=356 and cc>=146 and cc<150) then grbp<="110";
	end if;
	if (cc=187 and ll=356) then grbp<="110";
	end if;
	if (ll=356 and cc>=187 and cc<190) then grbp<="110";
	end if;
	if (cc=212 and ll=356) then grbp<="110";
	end if;
	if (cc=226 and ll=356) then grbp<="110";
	end if;
	if (ll=356 and cc>=226 and cc<228) then grbp<="110";
	end if;
	if (ll=357 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=357 and cc>=146 and cc<149) then grbp<="110";
	end if;
	if (cc=186 and ll=357) then grbp<="110";
	end if;
	if (cc=188 and ll=357) then grbp<="110";
	end if;
	if (ll=357 and cc>=188 and cc<192) then grbp<="110";
	end if;
	if (cc=226 and ll=357) then grbp<="110";
	end if;
	if (cc=18 and ll=358) then grbp<="110";
	end if;
	if (ll=358 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=358 and cc>=146 and cc<149) then grbp<="110";
	end if;
	if (ll=358 and cc>=186 and cc<188) then grbp<="110";
	end if;
	if (cc=192 and ll=358) then grbp<="110";
	end if;
	if (cc=211 and ll=358) then grbp<="110";
	end if;
	if (cc=225 and ll=358) then grbp<="110";
	end if;
	if (ll=358 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=359 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=359 and cc>=146 and cc<150) then grbp<="110";
	end if;
	if (ll=359 and cc>=185 and cc<188) then grbp<="110";
	end if;
	if (cc=225 and ll=359) then grbp<="110";
	end if;
	if (ll=359 and cc>=225 and cc<227) then grbp<="110";
	end if;
	if (ll=360 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=360 and cc>=146 and cc<152) then grbp<="110";
	end if;
	if (ll=360 and cc>=185 and cc<188) then grbp<="110";
	end if;
	if (cc=225 and ll=360) then grbp<="110";
	end if;
	if (cc=18 and ll=361) then grbp<="110";
	end if;
	if (ll=361 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=361 and cc>=147 and cc<150) then grbp<="110";
	end if;
	if (cc=187 and ll=361) then grbp<="110";
	end if;
	if (cc=192 and ll=361) then grbp<="110";
	end if;
	if (cc=224 and ll=361) then grbp<="110";
	end if;
	if (ll=361 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (ll=362 and cc>=18 and cc<20) then grbp<="110";
	end if;
	if (ll=362 and cc>=21 and cc<30) then grbp<="110";
	end if;
	if (ll=362 and cc>=145 and cc<152) then grbp<="110";
	end if;
	if (cc=187 and ll=362) then grbp<="110";
	end if;
	if (cc=210 and ll=362) then grbp<="110";
	end if;
	if (cc=224 and ll=362) then grbp<="110";
	end if;
	if (ll=362 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (ll=363 and cc>=18 and cc<24) then grbp<="110";
	end if;
	if (ll=363 and cc>=25 and cc<30) then grbp<="110";
	end if;
	if (ll=363 and cc>=145 and cc<151) then grbp<="110";
	end if;
	if (ll=363 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=210 and ll=363) then grbp<="110";
	end if;
	if (cc=224 and ll=363) then grbp<="110";
	end if;
	if (ll=363 and cc>=224 and cc<226) then grbp<="110";
	end if;
	if (ll=364 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=364 and cc>=147 and cc<151) then grbp<="110";
	end if;
	if (ll=364 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=210 and ll=364) then grbp<="110";
	end if;
	if (cc=224 and ll=364) then grbp<="110";
	end if;
	if (cc=18 and ll=365) then grbp<="110";
	end if;
	if (ll=365 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=365 and cc>=147 and cc<151) then grbp<="110";
	end if;
	if (cc=188 and ll=365) then grbp<="110";
	end if;
	if (ll=365 and cc>=188 and cc<190) then grbp<="110";
	end if;
	if (cc=223 and ll=365) then grbp<="110";
	end if;
	if (ll=365 and cc>=223 and cc<225) then grbp<="110";
	end if;
	if (ll=366 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=366 and cc>=146 and cc<152) then grbp<="110";
	end if;
	if (ll=366 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=223 and ll=366) then grbp<="110";
	end if;
	if (ll=366 and cc>=223 and cc<225) then grbp<="110";
	end if;
	if (ll=367 and cc>=18 and cc<22) then grbp<="110";
	end if;
	if (ll=367 and cc>=23 and cc<29) then grbp<="110";
	end if;
	if (cc=150 and ll=367) then grbp<="110";
	end if;
	if (ll=367 and cc>=150 and cc<153) then grbp<="110";
	end if;
	if (ll=367 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=223 and ll=367) then grbp<="110";
	end if;
	if (cc=18 and ll=368) then grbp<="110";
	end if;
	if (ll=368 and cc>=18 and cc<21) then grbp<="110";
	end if;
	if (ll=368 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (ll=368 and cc>=147 and cc<153) then grbp<="110";
	end if;
	if (ll=368 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=223 and ll=368) then grbp<="110";
	end if;
	if (cc=18 and ll=369) then grbp<="110";
	end if;
	if (ll=369 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=369 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (ll=369 and cc>=149 and cc<152) then grbp<="110";
	end if;
	if (ll=369 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=222 and ll=369) then grbp<="110";
	end if;
	if (ll=369 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=370 and cc>=18 and cc<23) then grbp<="110";
	end if;
	if (ll=370 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=370 and cc>=149 and cc<153) then grbp<="110";
	end if;
	if (ll=370 and cc>=185 and cc<189) then grbp<="110";
	end if;
	if (ll=370 and cc>=222 and cc<224) then grbp<="110";
	end if;
	if (ll=371 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=371 and cc>=148 and cc<154) then grbp<="110";
	end if;
	if (ll=371 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=222 and ll=371) then grbp<="110";
	end if;
	if (cc=18 and ll=372) then grbp<="110";
	end if;
	if (cc=20 and ll=372) then grbp<="110";
	end if;
	if (ll=372 and cc>=20 and cc<30) then grbp<="110";
	end if;
	if (ll=372 and cc>=148 and cc<154) then grbp<="110";
	end if;
	if (ll=372 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=222 and ll=372) then grbp<="110";
	end if;
	if (cc=18 and ll=373) then grbp<="110";
	end if;
	if (ll=373 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=373 and cc>=148 and cc<152) then grbp<="110";
	end if;
	if (cc=185 and ll=373) then grbp<="110";
	end if;
	if (ll=373 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (cc=210 and ll=373) then grbp<="110";
	end if;
	if (cc=221 and ll=373) then grbp<="110";
	end if;
	if (ll=373 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=374 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (cc=153 and ll=374) then grbp<="110";
	end if;
	if (ll=374 and cc>=153 and cc<155) then grbp<="110";
	end if;
	if (ll=374 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (ll=374 and cc>=210 and cc<212) then grbp<="110";
	end if;
	if (cc=221 and ll=374) then grbp<="110";
	end if;
	if (ll=374 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=375 and cc>=18 and cc<29) then grbp<="110";
	end if;
	if (ll=375 and cc>=148 and cc<152) then grbp<="110";
	end if;
	if (ll=375 and cc>=185 and cc<187) then grbp<="110";
	end if;
	if (ll=375 and cc>=211 and cc<216) then grbp<="110";
	end if;
	if (ll=375 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=376 and cc>=18 and cc<26) then grbp<="110";
	end if;
	if (ll=376 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (ll=376 and cc>=150 and cc<153) then grbp<="110";
	end if;
	if (ll=376 and cc>=154 and cc<156) then grbp<="110";
	end if;
	if (cc=187 and ll=376) then grbp<="110";
	end if;
	if (cc=190 and ll=376) then grbp<="110";
	end if;
	if (cc=193 and ll=376) then grbp<="110";
	end if;
	if (cc=211 and ll=376) then grbp<="110";
	end if;
	if (ll=376 and cc>=211 and cc<216) then grbp<="110";
	end if;
	if (ll=376 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=377 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=377 and cc>=150 and cc<156) then grbp<="110";
	end if;
	if (ll=377 and cc>=191 and cc<193) then grbp<="110";
	end if;
	if (ll=377 and cc>=212 and cc<215) then grbp<="110";
	end if;
	if (ll=377 and cc>=221 and cc<223) then grbp<="110";
	end if;
	if (ll=378 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (cc=150 and ll=378) then grbp<="110";
	end if;
	if (ll=378 and cc>=150 and cc<156) then grbp<="110";
	end if;
	if (ll=378 and cc>=192 and cc<195) then grbp<="110";
	end if;
	if (ll=378 and cc>=213 and cc<215) then grbp<="110";
	end if;
	if (cc=18 and ll=379) then grbp<="110";
	end if;
	if (ll=379 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (cc=151 and ll=379) then grbp<="110";
	end if;
	if (ll=379 and cc>=151 and cc<156) then grbp<="110";
	end if;
	if (ll=379 and cc>=194 and cc<196) then grbp<="110";
	end if;
	if (cc=214 and ll=379) then grbp<="110";
	end if;
	if (cc=221 and ll=379) then grbp<="110";
	end if;
	if (cc=18 and ll=380) then grbp<="110";
	end if;
	if (ll=380 and cc>=18 and cc<25) then grbp<="110";
	end if;
	if (ll=380 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (ll=380 and cc>=151 and cc<156) then grbp<="110";
	end if;
	if (cc=206 and ll=380) then grbp<="110";
	end if;
	if (ll=380 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (cc=220 and ll=380) then grbp<="110";
	end if;
	if (ll=380 and cc>=220 and cc<222) then grbp<="110";
	end if;
	if (ll=381 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=381 and cc>=152 and cc<154) then grbp<="110";
	end if;
	if (cc=207 and ll=381) then grbp<="110";
	end if;
	if (cc=214 and ll=381) then grbp<="110";
	end if;
	if (cc=220 and ll=381) then grbp<="110";
	end if;
	if (ll=381 and cc>=220 and cc<222) then grbp<="110";
	end if;
	if (ll=382 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=382 and cc>=152 and cc<157) then grbp<="110";
	end if;
	if (ll=382 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (cc=220 and ll=382) then grbp<="110";
	end if;
	if (ll=382 and cc>=220 and cc<222) then grbp<="110";
	end if;
	if (ll=383 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (cc=152 and ll=383) then grbp<="110";
	end if;
	if (ll=383 and cc>=152 and cc<158) then grbp<="110";
	end if;
	if (ll=383 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (cc=220 and ll=383) then grbp<="110";
	end if;
	if (cc=18 and ll=384) then grbp<="110";
	end if;
	if (ll=384 and cc>=18 and cc<30) then grbp<="110";
	end if;
	if (ll=384 and cc>=153 and cc<158) then grbp<="110";
	end if;
	if (ll=384 and cc>=204 and cc<208) then grbp<="110";
	end if;
	if (cc=219 and ll=384) then grbp<="110";
	end if;
	if (ll=384 and cc>=219 and cc<221) then grbp<="110";
	end if;
	if (ll=385 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=385 and cc>=151 and cc<157) then grbp<="110";
	end if;
	if (cc=205 and ll=385) then grbp<="110";
	end if;
	if (ll=385 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (cc=219 and ll=385) then grbp<="110";
	end if;
	if (ll=385 and cc>=219 and cc<221) then grbp<="110";
	end if;
	if (ll=386 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (ll=386 and cc>=23 and cc<30) then grbp<="110";
	end if;
	if (ll=386 and cc>=151 and cc<158) then grbp<="110";
	end if;
	if (ll=386 and cc>=205 and cc<208) then grbp<="110";
	end if;
	if (cc=219 and ll=386) then grbp<="110";
	end if;
	if (ll=386 and cc>=219 and cc<221) then grbp<="110";
	end if;
	if (ll=387 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=387 and cc>=152 and cc<156) then grbp<="110";
	end if;
	if (cc=206 and ll=387) then grbp<="110";
	end if;
	if (ll=387 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (ll=387 and cc>=209 and cc<211) then grbp<="110";
	end if;
	if (cc=218 and ll=387) then grbp<="110";
	end if;
	if (ll=387 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=388 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=388 and cc>=153 and cc<159) then grbp<="110";
	end if;
	if (ll=388 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (ll=388 and cc>=209 and cc<214) then grbp<="110";
	end if;
	if (ll=388 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=389 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=389 and cc>=153 and cc<160) then grbp<="110";
	end if;
	if (ll=389 and cc>=208 and cc<214) then grbp<="110";
	end if;
	if (ll=389 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=390 and cc>=18 and cc<26) then grbp<="110";
	end if;
	if (ll=390 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (ll=390 and cc>=154 and cc<159) then grbp<="110";
	end if;
	if (ll=390 and cc>=208 and cc<211) then grbp<="110";
	end if;
	if (cc=218 and ll=390) then grbp<="110";
	end if;
	if (ll=390 and cc>=218 and cc<220) then grbp<="110";
	end if;
	if (ll=391 and cc>=18 and cc<27) then grbp<="110";
	end if;
	if (ll=391 and cc>=28 and cc<30) then grbp<="110";
	end if;
	if (ll=391 and cc>=154 and cc<159) then grbp<="110";
	end if;
	if (ll=391 and cc>=207 and cc<213) then grbp<="110";
	end if;
	if (cc=19 and ll=392) then grbp<="110";
	end if;
	if (ll=392 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=392 and cc>=153 and cc<160) then grbp<="110";
	end if;
	if (cc=209 and ll=392) then grbp<="110";
	end if;
	if (ll=392 and cc>=209 and cc<213) then grbp<="110";
	end if;
	if (ll=392 and cc>=217 and cc<219) then grbp<="110";
	end if;
	if (ll=393 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (cc=154 and ll=393) then grbp<="110";
	end if;
	if (ll=393 and cc>=154 and cc<160) then grbp<="110";
	end if;
	if (cc=210 and ll=393) then grbp<="110";
	end if;
	if (ll=393 and cc>=210 and cc<213) then grbp<="110";
	end if;
	if (ll=393 and cc>=217 and cc<219) then grbp<="110";
	end if;
	if (ll=394 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=394 and cc>=154 and cc<160) then grbp<="110";
	end if;
	if (cc=209 and ll=394) then grbp<="110";
	end if;
	if (ll=394 and cc>=209 and cc<211) then grbp<="110";
	end if;
	if (cc=217 and ll=394) then grbp<="110";
	end if;
	if (cc=19 and ll=395) then grbp<="110";
	end if;
	if (ll=395 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=395 and cc>=153 and cc<161) then grbp<="110";
	end if;
	if (cc=206 and ll=395) then grbp<="110";
	end if;
	if (cc=209 and ll=395) then grbp<="110";
	end if;
	if (ll=395 and cc>=209 and cc<213) then grbp<="110";
	end if;
	if (ll=395 and cc>=216 and cc<218) then grbp<="110";
	end if;
	if (ll=396 and cc>=19 and cc<26) then grbp<="110";
	end if;
	if (ll=396 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (ll=396 and cc>=154 and cc<156) then grbp<="110";
	end if;
	if (ll=396 and cc>=157 and cc<160) then grbp<="110";
	end if;
	if (cc=209 and ll=396) then grbp<="110";
	end if;
	if (ll=396 and cc>=209 and cc<213) then grbp<="110";
	end if;
	if (ll=396 and cc>=216 and cc<218) then grbp<="110";
	end if;
	if (ll=397 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (cc=157 and ll=397) then grbp<="110";
	end if;
	if (ll=397 and cc>=157 and cc<160) then grbp<="110";
	end if;
	if (ll=397 and cc>=206 and cc<213) then grbp<="110";
	end if;
	if (ll=397 and cc>=215 and cc<217) then grbp<="110";
	end if;
	if (ll=398 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=398 and cc>=156 and cc<162) then grbp<="110";
	end if;
	if (ll=398 and cc>=206 and cc<214) then grbp<="110";
	end if;
	if (ll=398 and cc>=215 and cc<217) then grbp<="110";
	end if;
	if (ll=399 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=399 and cc>=156 and cc<162) then grbp<="110";
	end if;
	if (ll=399 and cc>=206 and cc<208) then grbp<="110";
	end if;
	if (ll=399 and cc>=210 and cc<216) then grbp<="110";
	end if;
	if (ll=400 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=400 and cc>=156 and cc<159) then grbp<="110";
	end if;
	if (ll=400 and cc>=161 and cc<163) then grbp<="110";
	end if;
	if (cc=206 and ll=400) then grbp<="110";
	end if;
	if (cc=211 and ll=400) then grbp<="110";
	end if;
	if (ll=400 and cc>=211 and cc<215) then grbp<="110";
	end if;
	if (ll=401 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=401 and cc>=157 and cc<160) then grbp<="110";
	end if;
	if (cc=206 and ll=401) then grbp<="110";
	end if;
	if (cc=211 and ll=401) then grbp<="110";
	end if;
	if (ll=401 and cc>=211 and cc<214) then grbp<="110";
	end if;
	if (ll=402 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=402 and cc>=158 and cc<162) then grbp<="110";
	end if;
	if (cc=211 and ll=402) then grbp<="110";
	end if;
	if (ll=402 and cc>=211 and cc<213) then grbp<="110";
	end if;
	if (ll=403 and cc>=19 and cc<25) then grbp<="110";
	end if;
	if (ll=403 and cc>=26 and cc<30) then grbp<="110";
	end if;
	if (cc=154 and ll=403) then grbp<="110";
	end if;
	if (cc=159 and ll=403) then grbp<="110";
	end if;
	if (ll=403 and cc>=159 and cc<162) then grbp<="110";
	end if;
	if (cc=211 and ll=403) then grbp<="110";
	end if;
	if (ll=403 and cc>=211 and cc<213) then grbp<="110";
	end if;
	if (ll=404 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=404 and cc>=159 and cc<162) then grbp<="110";
	end if;
	if (cc=210 and ll=404) then grbp<="110";
	end if;
	if (ll=404 and cc>=210 and cc<212) then grbp<="110";
	end if;
	if (ll=405 and cc>=19 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=405) then grbp<="110";
	end if;
	if (ll=405 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (cc=159 and ll=405) then grbp<="110";
	end if;
	if (cc=161 and ll=405) then grbp<="110";
	end if;
	if (ll=405 and cc>=161 and cc<163) then grbp<="110";
	end if;
	if (cc=206 and ll=405) then grbp<="110";
	end if;
	if (cc=211 and ll=405) then grbp<="110";
	end if;
	if (cc=19 and ll=406) then grbp<="110";
	end if;
	if (ll=406 and cc>=19 and cc<25) then grbp<="110";
	end if;
	if (ll=406 and cc>=26 and cc<30) then grbp<="110";
	end if;
	if (cc=150 and ll=406) then grbp<="110";
	end if;
	if (ll=406 and cc>=150 and cc<152) then grbp<="110";
	end if;
	if (cc=159 and ll=406) then grbp<="110";
	end if;
	if (cc=210 and ll=406) then grbp<="110";
	end if;
	if (ll=406 and cc>=210 and cc<212) then grbp<="110";
	end if;
	if (ll=407 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (cc=159 and ll=407) then grbp<="110";
	end if;
	if (cc=208 and ll=407) then grbp<="110";
	end if;
	if (cc=19 and ll=408) then grbp<="110";
	end if;
	if (ll=408 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (cc=159 and ll=408) then grbp<="110";
	end if;
	if (cc=161 and ll=408) then grbp<="110";
	end if;
	if (ll=408 and cc>=161 and cc<163) then grbp<="110";
	end if;
	if (cc=208 and ll=408) then grbp<="110";
	end if;
	if (ll=408 and cc>=208 and cc<210) then grbp<="110";
	end if;
	if (ll=409 and cc>=19 and cc<23) then grbp<="110";
	end if;
	if (ll=409 and cc>=24 and cc<26) then grbp<="110";
	end if;
	if (ll=409 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (cc=159 and ll=409) then grbp<="110";
	end if;
	if (cc=161 and ll=409) then grbp<="110";
	end if;
	if (ll=409 and cc>=161 and cc<163) then grbp<="110";
	end if;
	if (cc=207 and ll=409) then grbp<="110";
	end if;
	if (cc=19 and ll=410) then grbp<="110";
	end if;
	if (ll=410 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (ll=410 and cc>=23 and cc<26) then grbp<="110";
	end if;
	if (ll=410 and cc>=27 and cc<31) then grbp<="110";
	end if;
	if (cc=159 and ll=410) then grbp<="110";
	end if;
	if (cc=161 and ll=410) then grbp<="110";
	end if;
	if (cc=13 and ll=411) then grbp<="110";
	end if;
	if (cc=19 and ll=411) then grbp<="110";
	end if;
	if (ll=411 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (ll=411 and cc>=23 and cc<30) then grbp<="110";
	end if;
	if (ll=411 and cc>=151 and cc<153) then grbp<="110";
	end if;
	if (cc=159 and ll=411) then grbp<="110";
	end if;
	if (cc=161 and ll=411) then grbp<="110";
	end if;
	if (cc=19 and ll=412) then grbp<="110";
	end if;
	if (ll=412 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (cc=27 and ll=412) then grbp<="110";
	end if;
	if (ll=412 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (cc=159 and ll=412) then grbp<="110";
	end if;
	if (cc=19 and ll=413) then grbp<="110";
	end if;
	if (ll=413 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (cc=27 and ll=413) then grbp<="110";
	end if;
	if (ll=413 and cc>=27 and cc<30) then grbp<="110";
	end if;
	if (cc=146 and ll=413) then grbp<="110";
	end if;
	if (cc=154 and ll=413) then grbp<="110";
	end if;
	if (cc=163 and ll=413) then grbp<="110";
	end if;
	if (cc=19 and ll=414) then grbp<="110";
	end if;
	if (ll=414 and cc>=19 and cc<25) then grbp<="110";
	end if;
	if (ll=414 and cc>=26 and cc<30) then grbp<="110";
	end if;
	if (ll=414 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=414) then grbp<="110";
	end if;
	if (cc=19 and ll=415) then grbp<="110";
	end if;
	if (ll=415 and cc>=19 and cc<23) then grbp<="110";
	end if;
	if (ll=415 and cc>=26 and cc<29) then grbp<="110";
	end if;
	if (ll=415 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=415) then grbp<="110";
	end if;
	if (cc=19 and ll=416) then grbp<="110";
	end if;
	if (ll=416 and cc>=19 and cc<23) then grbp<="110";
	end if;
	if (cc=28 and ll=416) then grbp<="110";
	end if;
	if (cc=160 and ll=416) then grbp<="110";
	end if;
	if (ll=416 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=416) then grbp<="110";
	end if;
	if (cc=19 and ll=417) then grbp<="110";
	end if;
	if (ll=417 and cc>=19 and cc<23) then grbp<="110";
	end if;
	if (ll=417 and cc>=24 and cc<29) then grbp<="110";
	end if;
	if (ll=417 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=417) then grbp<="110";
	end if;
	if (cc=19 and ll=418) then grbp<="110";
	end if;
	if (ll=418 and cc>=19 and cc<30) then grbp<="110";
	end if;
	if (ll=418 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=418) then grbp<="110";
	end if;
	if (cc=19 and ll=419) then grbp<="110";
	end if;
	if (ll=419 and cc>=19 and cc<29) then grbp<="110";
	end if;
	if (cc=160 and ll=419) then grbp<="110";
	end if;
	if (cc=162 and ll=419) then grbp<="110";
	end if;
	if (ll=419 and cc>=162 and cc<164) then grbp<="110";
	end if;
	if (cc=19 and ll=420) then grbp<="110";
	end if;
	if (ll=420 and cc>=19 and cc<29) then grbp<="110";
	end if;
	if (cc=160 and ll=420) then grbp<="110";
	end if;
	if (ll=420 and cc>=160 and cc<162) then grbp<="110";
	end if;
	if (ll=421 and cc>=19 and cc<29) then grbp<="110";
	end if;
	if (ll=421 and cc>=160 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=421) then grbp<="110";
	end if;
	if (ll=421 and cc>=163 and cc<165) then grbp<="110";
	end if;
	if (ll=422 and cc>=19 and cc<24) then grbp<="110";
	end if;
	if (cc=27 and ll=422) then grbp<="110";
	end if;
	if (ll=422 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=159 and ll=422) then grbp<="110";
	end if;
	if (ll=422 and cc>=159 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=422) then grbp<="110";
	end if;
	if (cc=19 and ll=423) then grbp<="110";
	end if;
	if (ll=423 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (cc=25 and ll=423) then grbp<="110";
	end if;
	if (cc=27 and ll=423) then grbp<="110";
	end if;
	if (ll=423 and cc>=27 and cc<29) then grbp<="110";
	end if;
	if (cc=159 and ll=423) then grbp<="110";
	end if;
	if (ll=423 and cc>=159 and cc<163) then grbp<="110";
	end if;
	if (cc=163 and ll=423) then grbp<="110";
	end if;
	if (cc=19 and ll=424) then grbp<="110";
	end if;
	if (ll=424 and cc>=19 and cc<22) then grbp<="110";
	end if;
	if (ll=424 and cc>=23 and cc<26) then grbp<="110";
	end if;
	if (cc=157 and ll=424) then grbp<="110";
	end if;
	if (cc=159 and ll=424) then grbp<="110";
	end if;
	if (ll=424 and cc>=159 and cc<163) then grbp<="110";
	end if;

	if (cc=129 and ll=148) then grbp<="001";
	end if;
	if (cc=140 and ll=151) then grbp<="001";
	end if;
	if (cc=132 and ll=153) then grbp<="001";
	end if;
	if (cc=128 and ll=157) then grbp<="001";
	end if;
	if (cc=128 and ll=158) then grbp<="001";
	end if;
	if (cc=132 and ll=160) then grbp<="001";
	end if;
	if (cc=131 and ll=161) then grbp<="001";
	end if;
	if (cc=131 and ll=162) then grbp<="001";
	end if;
	if (cc=128 and ll=164) then grbp<="001";
	end if;
	if (cc=127 and ll=166) then grbp<="001";
	end if;
	if (ll=167 and cc>=127 and cc<129) then grbp<="001";
	end if;
	if (cc=126 and ll=170) then grbp<="001";
	end if;
	if (cc=126 and ll=176) then grbp<="001";
	end if;
	if (ll=178 and cc>=126 and cc<128) then grbp<="001";
	end if;
	if (cc=103 and ll=207) then grbp<="001";
	end if;
	if (cc=103 and ll=208) then grbp<="001";
	end if;
	if (cc=85 and ll=214) then grbp<="001";
	end if;
	if (cc=71 and ll=217) then grbp<="001";
	end if;
	if (cc=70 and ll=219) then grbp<="001";
	end if;
	if (cc=64 and ll=228) then grbp<="001";
	end if;
	if (cc=72 and ll=229) then grbp<="001";
	end if;
	if (cc=77 and ll=229) then grbp<="001";
	end if;
	if (cc=72 and ll=230) then grbp<="001";
	end if;
	if (cc=72 and ll=231) then grbp<="001";
	end if;
	if (cc=77 and ll=231) then grbp<="001";
	end if;
	if (cc=65 and ll=232) then grbp<="001";
	end if;
	if (cc=75 and ll=240) then grbp<="001";
	end if;
	if (ll=241 and cc>=75 and cc<77) then grbp<="001";
	end if;
	if (cc=59 and ll=247) then grbp<="001";
	end if;
	if (cc=61 and ll=248) then grbp<="001";
	end if;
	if (cc=64 and ll=248) then grbp<="001";
	end if;
	if (cc=60 and ll=251) then grbp<="001";
	end if;
	if (cc=60 and ll=252) then grbp<="001";
	end if;
	if (cc=57 and ll=255) then grbp<="001";
	end if;
	if (cc=59 and ll=255) then grbp<="001";
	end if;
	if (cc=55 and ll=256) then grbp<="001";
	end if;
	if (ll=258 and cc>=55 and cc<57) then grbp<="001";
	end if;
	if (cc=51 and ll=260) then grbp<="001";
	end if;
	if (cc=53 and ll=260) then grbp<="001";
	end if;
	if (cc=64 and ll=260) then grbp<="001";
	end if;
	if (cc=60 and ll=267) then grbp<="001";
	end if;
	if (ll=268 and cc>=60 and cc<62) then grbp<="001";
	end if;
	if (cc=60 and ll=269) then grbp<="001";
	end if;
	if (ll=269 and cc>=60 and cc<62) then grbp<="001";
	end if;
	if (cc=59 and ll=270) then grbp<="001";
	end if;
	if (cc=52 and ll=271) then grbp<="001";
	end if;
	if (cc=59 and ll=273) then grbp<="001";
	end if;
	if (cc=59 and ll=278) then grbp<="001";
	end if;
	if (cc=64 and ll=281) then grbp<="001";
	end if;
	if (cc=68 and ll=288) then grbp<="001";
	end if;
	if (cc=68 and ll=289) then grbp<="001";
	end if;
	if (cc=56 and ll=290) then grbp<="001";
	end if;
	if (cc=56 and ll=291) then grbp<="001";
	end if;
	if (cc=60 and ll=294) then grbp<="001";
	end if;
	if (ll=294 and cc>=60 and cc<63) then grbp<="001";
	end if;
	if (cc=54 and ll=297) then grbp<="001";
	end if;
	if (cc=54 and ll=298) then grbp<="001";
	end if;
	if (cc=62 and ll=299) then grbp<="001";
	end if;
	if (cc=60 and ll=301) then grbp<="001";
	end if;
	if (cc=50 and ll=302) then grbp<="001";
	end if;
	if (cc=54 and ll=302) then grbp<="001";
	end if;
	if (cc=54 and ll=303) then grbp<="001";
	end if;
	if (cc=59 and ll=303) then grbp<="001";
	end if;
	if (cc=66 and ll=303) then grbp<="001";
	end if;
	if (cc=64 and ll=305) then grbp<="001";
	end if;
	if (cc=67 and ll=306) then grbp<="001";
	end if;
	if (cc=60 and ll=307) then grbp<="001";
	end if;
	if (cc=58 and ll=308) then grbp<="001";
	end if;
	if (cc=65 and ll=309) then grbp<="001";
	end if;
	if (cc=58 and ll=310) then grbp<="001";
	end if;
	if (cc=67 and ll=312) then grbp<="001";
	end if;
	if (cc=62 and ll=315) then grbp<="001";
	end if;
	if (cc=64 and ll=318) then grbp<="001";
	end if;
	if (cc=55 and ll=319) then grbp<="001";
	end if;
	if (cc=69 and ll=322) then grbp<="001";
	end if;
	if (cc=66 and ll=325) then grbp<="001";
	end if;
	if (cc=69 and ll=325) then grbp<="001";
	end if;
	if (cc=69 and ll=326) then grbp<="001";
	end if;
	if (ll=327 and cc>=69 and cc<71) then grbp<="001";
	end if;
	if (ll=328 and cc>=62 and cc<65) then grbp<="001";
	end if;
	if (cc=72 and ll=328) then grbp<="001";
	end if;
	if (cc=69 and ll=329) then grbp<="001";
	end if;
	if (cc=72 and ll=329) then grbp<="001";
	end if;
	if (cc=68 and ll=331) then grbp<="001";
	end if;
	if (ll=331 and cc>=68 and cc<70) then grbp<="001";
	end if;
	if (cc=69 and ll=332) then grbp<="001";
	end if;
	if (ll=332 and cc>=69 and cc<71) then grbp<="001";
	end if;
	if (ll=345 and cc>=68 and cc<70) then grbp<="001";
	end if;
	if (cc=71 and ll=347) then grbp<="001";
	end if;
	if (ll=348 and cc>=71 and cc<73) then grbp<="001";
	end if;
	if (cc=68 and ll=354) then grbp<="001";
	end if;
	if (cc=68 and ll=357) then grbp<="001";
	end if;
	if (cc=72 and ll=357) then grbp<="001";
	end if;
	if (cc=75 and ll=357) then grbp<="001";
	end if;
	if (cc=75 and ll=358) then grbp<="001";
	end if;
	if (cc=49 and ll=359) then grbp<="001";
	end if;
	if (cc=75 and ll=362) then grbp<="001";
	end if;
	if (cc=70 and ll=363) then grbp<="001";
	end if;
	if (cc=74 and ll=363) then grbp<="001";
	end if;
	if (ll=363 and cc>=74 and cc<76) then grbp<="001";
	end if;
	if (cc=87 and ll=366) then grbp<="001";
	end if;
	if (cc=73 and ll=368) then grbp<="001";
	end if;
	if (cc=73 and ll=369) then grbp<="001";
	end if;
	if (cc=73 and ll=371) then grbp<="001";
	end if;
	if (cc=75 and ll=371) then grbp<="001";
	end if;
	if (cc=73 and ll=372) then grbp<="001";
	end if;
	if (cc=71 and ll=373) then grbp<="001";
	end if;
	if (cc=73 and ll=373) then grbp<="001";
	end if;
	if (cc=78 and ll=374) then grbp<="001";
	end if;
	if (cc=74 and ll=375) then grbp<="001";
	end if;
	if (cc=78 and ll=375) then grbp<="001";
	end if;
	if (cc=81 and ll=377) then grbp<="001";
	end if;
	if (cc=70 and ll=378) then grbp<="001";
	end if;
	if (cc=68 and ll=385) then grbp<="001";
	end if;
	if (ll=394 and cc>=68 and cc<71) then grbp<="001";
	end if;
	if (cc=76 and ll=400) then grbp<="001";
	end if;
	if (cc=75 and ll=406) then grbp<="001";
	end if;
	if (cc=78 and ll=412) then grbp<="001";
	end if;
	if (cc=80 and ll=419) then grbp<="001";
	end if;

	if (cc=104 and ll=39) then grbp<="011";
	end if;
	if (cc=100 and ll=40) then grbp<="011";
	end if;
	if (ll=40 and cc>=100 and cc<105) then grbp<="011";
	end if;
	if (cc=97 and ll=41) then grbp<="011";
	end if;
	if (ll=41 and cc>=97 and cc<99) then grbp<="011";
	end if;
	if (ll=41 and cc>=102 and cc<104) then grbp<="011";
	end if;
	if (ll=42 and cc>=95 and cc<97) then grbp<="011";
	end if;
	if (cc=100 and ll=42) then grbp<="011";
	end if;
	if (cc=93 and ll=43) then grbp<="011";
	end if;
	if (ll=43 and cc>=93 and cc<96) then grbp<="011";
	end if;
	if (cc=102 and ll=43) then grbp<="011";
	end if;
	if (cc=126 and ll=43) then grbp<="011";
	end if;
	if (cc=96 and ll=44) then grbp<="011";
	end if;
	if (cc=102 and ll=44) then grbp<="011";
	end if;
	if (cc=93 and ll=45) then grbp<="011";
	end if;
	if (cc=95 and ll=45) then grbp<="011";
	end if;
	if (ll=45 and cc>=95 and cc<97) then grbp<="011";
	end if;
	if (cc=92 and ll=46) then grbp<="011";
	end if;
	if (ll=46 and cc>=92 and cc<94) then grbp<="011";
	end if;
	if (cc=98 and ll=46) then grbp<="011";
	end if;
	if (ll=46 and cc>=98 and cc<100) then grbp<="011";
	end if;
	if (ll=47 and cc>=86 and cc<88) then grbp<="011";
	end if;
	if (cc=96 and ll=47) then grbp<="011";
	end if;
	if (cc=102 and ll=47) then grbp<="011";
	end if;
	if (ll=47 and cc>=102 and cc<104) then grbp<="011";
	end if;
	if (ll=48 and cc>=83 and cc<87) then grbp<="011";
	end if;
	if (cc=104 and ll=48) then grbp<="011";
	end if;
	if (cc=131 and ll=48) then grbp<="011";
	end if;
	if (cc=81 and ll=49) then grbp<="011";
	end if;
	if (cc=84 and ll=49) then grbp<="011";
	end if;
	if (ll=49 and cc>=84 and cc<86) then grbp<="011";
	end if;
	if (cc=102 and ll=49) then grbp<="011";
	end if;
	if (cc=82 and ll=50) then grbp<="011";
	end if;
	if (cc=101 and ll=51) then grbp<="011";
	end if;
	if (cc=105 and ll=51) then grbp<="011";
	end if;
	if (cc=103 and ll=53) then grbp<="011";
	end if;
	if (cc=109 and ll=53) then grbp<="011";
	end if;
	if (cc=104 and ll=54) then grbp<="011";
	end if;
	if (cc=108 and ll=54) then grbp<="011";
	end if;
	if (cc=102 and ll=55) then grbp<="011";
	end if;
	if (cc=104 and ll=55) then grbp<="011";
	end if;
	if (cc=107 and ll=55) then grbp<="011";
	end if;
	if (cc=104 and ll=56) then grbp<="011";
	end if;
	if (ll=58 and cc>=104 and cc<106) then grbp<="011";
	end if;
	if (cc=112 and ll=75) then grbp<="011";
	end if;
	if (cc=245 and ll=76) then grbp<="011";
	end if;
	if (cc=118 and ll=78) then grbp<="011";
	end if;
	if (cc=244 and ll=78) then grbp<="011";
	end if;
	if (cc=117 and ll=79) then grbp<="011";
	end if;
	if (cc=116 and ll=80) then grbp<="011";
	end if;
	if (cc=242 and ll=82) then grbp<="011";
	end if;
	if (cc=113 and ll=84) then grbp<="011";
	end if;
	if (cc=239 and ll=85) then grbp<="011";
	end if;
	if (cc=239 and ll=87) then grbp<="011";
	end if;
	if (cc=243 and ll=88) then grbp<="011";
	end if;
	if (cc=108 and ll=90) then grbp<="011";
	end if;
	if (cc=235 and ll=92) then grbp<="011";
	end if;
	if (cc=193 and ll=93) then grbp<="011";
	end if;
	if (cc=192 and ll=94) then grbp<="011";
	end if;
	if (cc=104 and ll=95) then grbp<="011";
	end if;
	if (cc=233 and ll=97) then grbp<="011";
	end if;
	if (cc=189 and ll=98) then grbp<="011";
	end if;
	if (cc=233 and ll=98) then grbp<="011";
	end if;
	if (cc=204 and ll=99) then grbp<="011";
	end if;
	if (cc=232 and ll=99) then grbp<="011";
	end if;
	if (cc=231 and ll=101) then grbp<="011";
	end if;
	if (cc=186 and ll=102) then grbp<="011";
	end if;
	if (cc=231 and ll=102) then grbp<="011";
	end if;
	if (cc=98 and ll=103) then grbp<="011";
	end if;
	if (cc=162 and ll=103) then grbp<="011";
	end if;
	if (cc=231 and ll=103) then grbp<="011";
	end if;
	if (cc=97 and ll=105) then grbp<="011";
	end if;
	if (cc=230 and ll=105) then grbp<="011";
	end if;
	if (cc=163 and ll=106) then grbp<="011";
	end if;
	if (cc=183 and ll=106) then grbp<="011";
	end if;
	if (cc=230 and ll=106) then grbp<="011";
	end if;
	if (cc=182 and ll=107) then grbp<="011";
	end if;
	if (cc=229 and ll=108) then grbp<="011";
	end if;
	if (cc=229 and ll=109) then grbp<="011";
	end if;
	if (cc=231 and ll=109) then grbp<="011";
	end if;
	if (ll=109 and cc>=231 and cc<233) then grbp<="011";
	end if;
	if (cc=103 and ll=111) then grbp<="011";
	end if;
	if (cc=228 and ll=111) then grbp<="011";
	end if;
	if (cc=231 and ll=111) then grbp<="011";
	end if;
	if (cc=103 and ll=112) then grbp<="011";
	end if;
	if (cc=177 and ll=112) then grbp<="011";
	end if;
	if (cc=232 and ll=113) then grbp<="011";
	end if;
	if (cc=89 and ll=117) then grbp<="011";
	end if;
	if (cc=118 and ll=117) then grbp<="011";
	end if;
	if (cc=90 and ll=120) then grbp<="011";
	end if;
	if (cc=87 and ll=121) then grbp<="011";
	end if;
	if (cc=229 and ll=121) then grbp<="011";
	end if;
	if (cc=224 and ll=122) then grbp<="011";
	end if;
	if (cc=100 and ll=123) then grbp<="011";
	end if;
	if (cc=114 and ll=123) then grbp<="011";
	end if;
	if (cc=223 and ll=124) then grbp<="011";
	end if;
	if (cc=87 and ll=125) then grbp<="011";
	end if;
	if (cc=228 and ll=125) then grbp<="011";
	end if;
	if (cc=98 and ll=126) then grbp<="011";
	end if;
	if (ll=128 and cc>=98 and cc<100) then grbp<="011";
	end if;
	if (cc=110 and ll=128) then grbp<="011";
	end if;
	if (cc=222 and ll=128) then grbp<="011";
	end if;
	if (cc=89 and ll=129) then grbp<="011";
	end if;
	if (cc=109 and ll=129) then grbp<="011";
	end if;
	if (cc=101 and ll=130) then grbp<="011";
	end if;
	if (cc=226 and ll=130) then grbp<="011";
	end if;
	if (cc=98 and ll=132) then grbp<="011";
	end if;
	if (cc=105 and ll=132) then grbp<="011";
	end if;
	if (cc=131 and ll=132) then grbp<="011";
	end if;
	if (cc=197 and ll=132) then grbp<="011";
	end if;
	if (cc=221 and ll=132) then grbp<="011";
	end if;
	if (cc=109 and ll=133) then grbp<="011";
	end if;
	if (cc=155 and ll=133) then grbp<="011";
	end if;
	if (cc=101 and ll=134) then grbp<="011";
	end if;
	if (ll=135 and cc>=101 and cc<103) then grbp<="011";
	end if;
	if (ll=136 and cc>=104 and cc<106) then grbp<="011";
	end if;
	if (cc=111 and ll=136) then grbp<="011";
	end if;
	if (cc=117 and ll=136) then grbp<="011";
	end if;
	if (cc=127 and ll=136) then grbp<="011";
	end if;
	if (cc=152 and ll=136) then grbp<="011";
	end if;
	if (cc=112 and ll=137) then grbp<="011";
	end if;
	if (cc=117 and ll=137) then grbp<="011";
	end if;
	if (cc=150 and ll=137) then grbp<="011";
	end if;
	if (cc=197 and ll=137) then grbp<="011";
	end if;
	if (cc=219 and ll=137) then grbp<="011";
	end if;
	if (cc=224 and ll=137) then grbp<="011";
	end if;
	if (cc=101 and ll=138) then grbp<="011";
	end if;
	if (cc=110 and ll=138) then grbp<="011";
	end if;
	if (cc=115 and ll=138) then grbp<="011";
	end if;
	if (ll=138 and cc>=115 and cc<118) then grbp<="011";
	end if;
	if (cc=150 and ll=138) then grbp<="011";
	end if;
	if (cc=197 and ll=138) then grbp<="011";
	end if;
	if (cc=220 and ll=138) then grbp<="011";
	end if;
	if (cc=110 and ll=139) then grbp<="011";
	end if;
	if (cc=113 and ll=139) then grbp<="011";
	end if;
	if (cc=116 and ll=139) then grbp<="011";
	end if;
	if (ll=139 and cc>=116 and cc<119) then grbp<="011";
	end if;
	if (cc=192 and ll=139) then grbp<="011";
	end if;
	if (cc=220 and ll=139) then grbp<="011";
	end if;
	if (cc=110 and ll=140) then grbp<="011";
	end if;
	if (ll=140 and cc>=110 and cc<112) then grbp<="011";
	end if;
	if (ll=140 and cc>=115 and cc<118) then grbp<="011";
	end if;
	if (cc=145 and ll=140) then grbp<="011";
	end if;
	if (cc=148 and ll=140) then grbp<="011";
	end if;
	if (cc=188 and ll=140) then grbp<="011";
	end if;
	if (cc=107 and ll=141) then grbp<="011";
	end if;
	if (cc=109 and ll=141) then grbp<="011";
	end if;
	if (cc=111 and ll=141) then grbp<="011";
	end if;
	if (ll=141 and cc>=111 and cc<113) then grbp<="011";
	end if;
	if (ll=141 and cc>=115 and cc<120) then grbp<="011";
	end if;
	if (cc=99 and ll=142) then grbp<="011";
	end if;
	if (cc=104 and ll=142) then grbp<="011";
	end if;
	if (cc=114 and ll=142) then grbp<="011";
	end if;
	if (cc=129 and ll=142) then grbp<="011";
	end if;
	if (cc=138 and ll=142) then grbp<="011";
	end if;
	if (cc=222 and ll=142) then grbp<="011";
	end if;
	if (cc=102 and ll=143) then grbp<="011";
	end if;
	if (cc=119 and ll=143) then grbp<="011";
	end if;
	if (cc=121 and ll=143) then grbp<="011";
	end if;
	if (cc=123 and ll=143) then grbp<="011";
	end if;
	if (cc=129 and ll=143) then grbp<="011";
	end if;
	if (ll=143 and cc>=129 and cc<134) then grbp<="011";
	end if;
	if (ll=143 and cc>=137 and cc<139) then grbp<="011";
	end if;
	if (cc=108 and ll=144) then grbp<="011";
	end if;
	if (cc=117 and ll=144) then grbp<="011";
	end if;
	if (cc=121 and ll=144) then grbp<="011";
	end if;
	if (ll=144 and cc>=121 and cc<123) then grbp<="011";
	end if;
	if (ll=144 and cc>=126 and cc<128) then grbp<="011";
	end if;
	if (ll=144 and cc>=132 and cc<134) then grbp<="011";
	end if;
	if (cc=138 and ll=144) then grbp<="011";
	end if;
	if (ll=144 and cc>=138 and cc<140) then grbp<="011";
	end if;
	if (cc=144 and ll=144) then grbp<="011";
	end if;
	if (ll=144 and cc>=144 and cc<146) then grbp<="011";
	end if;
	if (cc=108 and ll=145) then grbp<="011";
	end if;
	if (cc=117 and ll=145) then grbp<="011";
	end if;
	if (cc=122 and ll=145) then grbp<="011";
	end if;
	if (ll=145 and cc>=122 and cc<126) then grbp<="011";
	end if;
	if (cc=135 and ll=145) then grbp<="011";
	end if;
	if (cc=139 and ll=145) then grbp<="011";
	end if;
	if (ll=145 and cc>=139 and cc<141) then grbp<="011";
	end if;
	if (cc=219 and ll=145) then grbp<="011";
	end if;
	if (cc=101 and ll=146) then grbp<="011";
	end if;
	if (cc=104 and ll=146) then grbp<="011";
	end if;
	if (cc=106 and ll=146) then grbp<="011";
	end if;
	if (ll=146 and cc>=106 and cc<109) then grbp<="011";
	end if;
	if (cc=122 and ll=146) then grbp<="011";
	end if;
	if (ll=146 and cc>=122 and cc<128) then grbp<="011";
	end if;
	if (cc=133 and ll=146) then grbp<="011";
	end if;
	if (ll=146 and cc>=133 and cc<135) then grbp<="011";
	end if;
	if (cc=102 and ll=147) then grbp<="011";
	end if;
	if (cc=106 and ll=147) then grbp<="011";
	end if;
	if (cc=117 and ll=147) then grbp<="011";
	end if;
	if (cc=121 and ll=147) then grbp<="011";
	end if;
	if (ll=147 and cc>=121 and cc<128) then grbp<="011";
	end if;
	if (cc=216 and ll=147) then grbp<="011";
	end if;
	if (cc=102 and ll=148) then grbp<="011";
	end if;
	if (cc=105 and ll=148) then grbp<="011";
	end if;
	if (ll=148 and cc>=105 and cc<107) then grbp<="011";
	end if;
	if (ll=148 and cc>=117 and cc<119) then grbp<="011";
	end if;
	if (ll=148 and cc>=121 and cc<127) then grbp<="011";
	end if;
	if (cc=193 and ll=148) then grbp<="011";
	end if;
	if (cc=117 and ll=149) then grbp<="011";
	end if;
	if (ll=149 and cc>=117 and cc<119) then grbp<="011";
	end if;
	if (ll=149 and cc>=120 and cc<124) then grbp<="011";
	end if;
	if (cc=104 and ll=150) then grbp<="011";
	end if;
	if (cc=114 and ll=150) then grbp<="011";
	end if;
	if (cc=116 and ll=150) then grbp<="011";
	end if;
	if (ll=150 and cc>=116 and cc<122) then grbp<="011";
	end if;
	if (ll=150 and cc>=128 and cc<130) then grbp<="011";
	end if;
	if (cc=145 and ll=150) then grbp<="011";
	end if;
	if (cc=105 and ll=151) then grbp<="011";
	end if;
	if (cc=109 and ll=151) then grbp<="011";
	end if;
	if (cc=112 and ll=151) then grbp<="011";
	end if;
	if (ll=151 and cc>=112 and cc<115) then grbp<="011";
	end if;
	if (cc=120 and ll=151) then grbp<="011";
	end if;
	if (ll=151 and cc>=120 and cc<122) then grbp<="011";
	end if;
	if (ll=151 and cc>=127 and cc<129) then grbp<="011";
	end if;
	if (cc=106 and ll=152) then grbp<="011";
	end if;
	if (cc=111 and ll=152) then grbp<="011";
	end if;
	if (ll=152 and cc>=111 and cc<115) then grbp<="011";
	end if;
	if (ll=152 and cc>=119 and cc<121) then grbp<="011";
	end if;
	if (cc=140 and ll=152) then grbp<="011";
	end if;
	if (cc=144 and ll=152) then grbp<="011";
	end if;
	if (cc=219 and ll=152) then grbp<="011";
	end if;
	if (cc=110 and ll=153) then grbp<="011";
	end if;
	if (cc=119 and ll=153) then grbp<="011";
	end if;
	if (ll=153 and cc>=119 and cc<122) then grbp<="011";
	end if;
	if (ll=153 and cc>=125 and cc<127) then grbp<="011";
	end if;
	if (ll=154 and cc>=107 and cc<111) then grbp<="011";
	end if;
	if (ll=154 and cc>=119 and cc<126) then grbp<="011";
	end if;
	if (cc=132 and ll=154) then grbp<="011";
	end if;
	if (cc=139 and ll=154) then grbp<="011";
	end if;
	if (cc=106 and ll=155) then grbp<="011";
	end if;
	if (ll=155 and cc>=106 and cc<110) then grbp<="011";
	end if;
	if (ll=155 and cc>=118 and cc<121) then grbp<="011";
	end if;
	if (cc=124 and ll=155) then grbp<="011";
	end if;
	if (cc=126 and ll=155) then grbp<="011";
	end if;
	if (ll=155 and cc>=126 and cc<128) then grbp<="011";
	end if;
	if (cc=214 and ll=155) then grbp<="011";
	end if;
	if (cc=106 and ll=156) then grbp<="011";
	end if;
	if (cc=118 and ll=156) then grbp<="011";
	end if;
	if (cc=120 and ll=156) then grbp<="011";
	end if;
	if (cc=124 and ll=156) then grbp<="011";
	end if;
	if (cc=126 and ll=156) then grbp<="011";
	end if;
	if (cc=132 and ll=156) then grbp<="011";
	end if;
	if (cc=215 and ll=156) then grbp<="011";
	end if;
	if (cc=100 and ll=157) then grbp<="011";
	end if;
	if (cc=118 and ll=157) then grbp<="011";
	end if;
	if (ll=157 and cc>=118 and cc<120) then grbp<="011";
	end if;
	if (cc=137 and ll=157) then grbp<="011";
	end if;
	if (cc=174 and ll=157) then grbp<="011";
	end if;
	if (cc=100 and ll=158) then grbp<="011";
	end if;
	if (cc=109 and ll=158) then grbp<="011";
	end if;
	if (cc=117 and ll=158) then grbp<="011";
	end if;
	if (cc=119 and ll=158) then grbp<="011";
	end if;
	if (cc=125 and ll=158) then grbp<="011";
	end if;
	if (cc=174 and ll=158) then grbp<="011";
	end if;
	if (ll=158 and cc>=174 and cc<176) then grbp<="011";
	end if;
	if (cc=117 and ll=159) then grbp<="011";
	end if;
	if (ll=159 and cc>=117 and cc<120) then grbp<="011";
	end if;
	if (cc=127 and ll=159) then grbp<="011";
	end if;
	if (cc=174 and ll=159) then grbp<="011";
	end if;
	if (ll=159 and cc>=174 and cc<176) then grbp<="011";
	end if;
	if (cc=116 and ll=160) then grbp<="011";
	end if;
	if (ll=160 and cc>=116 and cc<119) then grbp<="011";
	end if;
	if (cc=174 and ll=160) then grbp<="011";
	end if;
	if (ll=160 and cc>=174 and cc<178) then grbp<="011";
	end if;
	if (cc=106 and ll=161) then grbp<="011";
	end if;
	if (cc=116 and ll=161) then grbp<="011";
	end if;
	if (cc=123 and ll=161) then grbp<="011";
	end if;
	if (cc=175 and ll=161) then grbp<="011";
	end if;
	if (ll=161 and cc>=175 and cc<177) then grbp<="011";
	end if;
	if (cc=116 and ll=162) then grbp<="011";
	end if;
	if (cc=123 and ll=162) then grbp<="011";
	end if;
	if (cc=175 and ll=162) then grbp<="011";
	end if;
	if (ll=162 and cc>=175 and cc<177) then grbp<="011";
	end if;
	if (ll=163 and cc>=115 and cc<117) then grbp<="011";
	end if;
	if (ll=163 and cc>=122 and cc<124) then grbp<="011";
	end if;
	if (cc=131 and ll=163) then grbp<="011";
	end if;
	if (cc=133 and ll=163) then grbp<="011";
	end if;
	if (cc=175 and ll=163) then grbp<="011";
	end if;
	if (ll=163 and cc>=175 and cc<177) then grbp<="011";
	end if;
	if (cc=115 and ll=164) then grbp<="011";
	end if;
	if (cc=121 and ll=164) then grbp<="011";
	end if;
	if (ll=164 and cc>=121 and cc<123) then grbp<="011";
	end if;
	if (ll=164 and cc>=124 and cc<126) then grbp<="011";
	end if;
	if (cc=171 and ll=164) then grbp<="011";
	end if;
	if (cc=175 and ll=164) then grbp<="011";
	end if;
	if (ll=164 and cc>=175 and cc<177) then grbp<="011";
	end if;
	if (cc=123 and ll=165) then grbp<="011";
	end if;
	if (ll=165 and cc>=123 and cc<125) then grbp<="011";
	end if;
	if (cc=176 and ll=165) then grbp<="011";
	end if;
	if (cc=109 and ll=166) then grbp<="011";
	end if;
	if (cc=114 and ll=166) then grbp<="011";
	end if;
	if (ll=166 and cc>=114 and cc<116) then grbp<="011";
	end if;
	if (cc=135 and ll=166) then grbp<="011";
	end if;
	if (cc=171 and ll=166) then grbp<="011";
	end if;
	if (ll=166 and cc>=171 and cc<173) then grbp<="011";
	end if;
	if (cc=176 and ll=166) then grbp<="011";
	end if;
	if (ll=166 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (cc=172 and ll=167) then grbp<="011";
	end if;
	if (cc=174 and ll=167) then grbp<="011";
	end if;
	if (cc=176 and ll=167) then grbp<="011";
	end if;
	if (ll=167 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (cc=130 and ll=168) then grbp<="011";
	end if;
	if (ll=168 and cc>=130 and cc<132) then grbp<="011";
	end if;
	if (cc=108 and ll=169) then grbp<="011";
	end if;
	if (cc=123 and ll=169) then grbp<="011";
	end if;
	if (cc=127 and ll=169) then grbp<="011";
	end if;
	if (cc=130 and ll=169) then grbp<="011";
	end if;
	if (cc=173 and ll=169) then grbp<="011";
	end if;
	if (cc=177 and ll=169) then grbp<="011";
	end if;
	if (ll=169 and cc>=177 and cc<179) then grbp<="011";
	end if;
	if (cc=108 and ll=170) then grbp<="011";
	end if;
	if (cc=123 and ll=170) then grbp<="011";
	end if;
	if (cc=127 and ll=170) then grbp<="011";
	end if;
	if (cc=129 and ll=170) then grbp<="011";
	end if;
	if (cc=173 and ll=170) then grbp<="011";
	end if;
	if (cc=177 and ll=170) then grbp<="011";
	end if;
	if (ll=170 and cc>=177 and cc<179) then grbp<="011";
	end if;
	if (ll=171 and cc>=83 and cc<86) then grbp<="011";
	end if;
	if (cc=108 and ll=171) then grbp<="011";
	end if;
	if (cc=123 and ll=171) then grbp<="011";
	end if;
	if (cc=126 and ll=171) then grbp<="011";
	end if;
	if (ll=171 and cc>=126 and cc<130) then grbp<="011";
	end if;
	if (cc=173 and ll=171) then grbp<="011";
	end if;
	if (ll=171 and cc>=173 and cc<176) then grbp<="011";
	end if;
	if (cc=214 and ll=171) then grbp<="011";
	end if;
	if (cc=83 and ll=172) then grbp<="011";
	end if;
	if (ll=172 and cc>=83 and cc<89) then grbp<="011";
	end if;
	if (cc=107 and ll=172) then grbp<="011";
	end if;
	if (ll=172 and cc>=107 and cc<109) then grbp<="011";
	end if;
	if (cc=126 and ll=172) then grbp<="011";
	end if;
	if (ll=172 and cc>=126 and cc<128) then grbp<="011";
	end if;
	if (cc=131 and ll=172) then grbp<="011";
	end if;
	if (cc=169 and ll=172) then grbp<="011";
	end if;
	if (cc=174 and ll=172) then grbp<="011";
	end if;
	if (ll=172 and cc>=174 and cc<176) then grbp<="011";
	end if;
	if (cc=86 and ll=173) then grbp<="011";
	end if;
	if (ll=173 and cc>=86 and cc<89) then grbp<="011";
	end if;
	if (ll=173 and cc>=90 and cc<92) then grbp<="011";
	end if;
	if (ll=173 and cc>=107 and cc<109) then grbp<="011";
	end if;
	if (cc=126 and ll=173) then grbp<="011";
	end if;
	if (ll=173 and cc>=126 and cc<130) then grbp<="011";
	end if;
	if (cc=174 and ll=173) then grbp<="011";
	end if;
	if (ll=173 and cc>=174 and cc<178) then grbp<="011";
	end if;
	if (ll=174 and cc>=87 and cc<90) then grbp<="011";
	end if;
	if (cc=128 and ll=174) then grbp<="011";
	end if;
	if (ll=174 and cc>=128 and cc<131) then grbp<="011";
	end if;
	if (ll=174 and cc>=174 and cc<178) then grbp<="011";
	end if;
	if (cc=128 and ll=175) then grbp<="011";
	end if;
	if (ll=175 and cc>=128 and cc<130) then grbp<="011";
	end if;
	if (cc=175 and ll=175) then grbp<="011";
	end if;
	if (ll=175 and cc>=175 and cc<178) then grbp<="011";
	end if;
	if (ll=176 and cc>=128 and cc<131) then grbp<="011";
	end if;
	if (ll=176 and cc>=175 and cc<178) then grbp<="011";
	end if;
	if (cc=128 and ll=177) then grbp<="011";
	end if;
	if (ll=177 and cc>=128 and cc<130) then grbp<="011";
	end if;
	if (ll=177 and cc>=175 and cc<178) then grbp<="011";
	end if;
	if (ll=178 and cc>=108 and cc<110) then grbp<="011";
	end if;
	if (cc=129 and ll=178) then grbp<="011";
	end if;
	if (cc=175 and ll=178) then grbp<="011";
	end if;
	if (ll=178 and cc>=175 and cc<178) then grbp<="011";
	end if;
	if (cc=109 and ll=179) then grbp<="011";
	end if;
	if (cc=123 and ll=179) then grbp<="011";
	end if;
	if (cc=127 and ll=179) then grbp<="011";
	end if;
	if (cc=176 and ll=179) then grbp<="011";
	end if;
	if (ll=179 and cc>=176 and cc<179) then grbp<="011";
	end if;
	if (ll=180 and cc>=109 and cc<111) then grbp<="011";
	end if;
	if (ll=180 and cc>=126 and cc<128) then grbp<="011";
	end if;
	if (ll=180 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (cc=109 and ll=181) then grbp<="011";
	end if;
	if (ll=181 and cc>=109 and cc<112) then grbp<="011";
	end if;
	if (cc=176 and ll=181) then grbp<="011";
	end if;
	if (ll=181 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (cc=110 and ll=182) then grbp<="011";
	end if;
	if (ll=182 and cc>=110 and cc<112) then grbp<="011";
	end if;
	if (cc=127 and ll=182) then grbp<="011";
	end if;
	if (cc=176 and ll=182) then grbp<="011";
	end if;
	if (ll=182 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (ll=183 and cc>=110 and cc<112) then grbp<="011";
	end if;
	if (ll=183 and cc>=127 and cc<129) then grbp<="011";
	end if;
	if (ll=183 and cc>=176 and cc<178) then grbp<="011";
	end if;
	if (cc=127 and ll=184) then grbp<="011";
	end if;
	if (ll=184 and cc>=127 and cc<129) then grbp<="011";
	end if;
	if (cc=111 and ll=185) then grbp<="011";
	end if;
	if (cc=123 and ll=185) then grbp<="011";
	end if;
	if (cc=127 and ll=185) then grbp<="011";
	end if;
	if (ll=185 and cc>=127 and cc<129) then grbp<="011";
	end if;
	if (cc=128 and ll=186) then grbp<="011";
	end if;
	if (cc=111 and ll=187) then grbp<="011";
	end if;
	if (cc=122 and ll=187) then grbp<="011";
	end if;
	if (cc=128 and ll=187) then grbp<="011";
	end if;
	if (cc=143 and ll=187) then grbp<="011";
	end if;
	if (cc=90 and ll=188) then grbp<="011";
	end if;
	if (cc=108 and ll=188) then grbp<="011";
	end if;
	if (cc=111 and ll=188) then grbp<="011";
	end if;
	if (cc=128 and ll=188) then grbp<="011";
	end if;
	if (cc=177 and ll=188) then grbp<="011";
	end if;
	if (cc=107 and ll=189) then grbp<="011";
	end if;
	if (ll=189 and cc>=107 and cc<109) then grbp<="011";
	end if;
	if (cc=177 and ll=189) then grbp<="011";
	end if;
	if (cc=108 and ll=190) then grbp<="011";
	end if;
	if (cc=112 and ll=190) then grbp<="011";
	end if;
	if (cc=128 and ll=190) then grbp<="011";
	end if;
	if (cc=141 and ll=190) then grbp<="011";
	end if;
	if (cc=177 and ll=190) then grbp<="011";
	end if;
	if (cc=109 and ll=191) then grbp<="011";
	end if;
	if (cc=111 and ll=191) then grbp<="011";
	end if;
	if (ll=191 and cc>=111 and cc<113) then grbp<="011";
	end if;
	if (cc=107 and ll=192) then grbp<="011";
	end if;
	if (cc=112 and ll=192) then grbp<="011";
	end if;
	if (cc=140 and ll=192) then grbp<="011";
	end if;
	if (cc=106 and ll=193) then grbp<="011";
	end if;
	if (cc=112 and ll=193) then grbp<="011";
	end if;
	if (cc=84 and ll=194) then grbp<="011";
	end if;
	if (ll=194 and cc>=84 and cc<86) then grbp<="011";
	end if;
	if (cc=128 and ll=194) then grbp<="011";
	end if;
	if (cc=85 and ll=195) then grbp<="011";
	end if;
	if (cc=112 and ll=195) then grbp<="011";
	end if;
	if (ll=195 and cc>=112 and cc<114) then grbp<="011";
	end if;
	if (cc=137 and ll=195) then grbp<="011";
	end if;
	if (cc=228 and ll=195) then grbp<="011";
	end if;
	if (cc=75 and ll=196) then grbp<="011";
	end if;
	if (ll=196 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (cc=113 and ll=196) then grbp<="011";
	end if;
	if (cc=128 and ll=196) then grbp<="011";
	end if;
	if (cc=136 and ll=196) then grbp<="011";
	end if;
	if (cc=138 and ll=196) then grbp<="011";
	end if;
	if (cc=178 and ll=196) then grbp<="011";
	end if;
	if (cc=237 and ll=196) then grbp<="011";
	end if;
	if (cc=74 and ll=197) then grbp<="011";
	end if;
	if (ll=197 and cc>=74 and cc<77) then grbp<="011";
	end if;
	if (cc=236 and ll=197) then grbp<="011";
	end if;
	if (cc=73 and ll=198) then grbp<="011";
	end if;
	if (ll=198 and cc>=73 and cc<77) then grbp<="011";
	end if;
	if (cc=108 and ll=198) then grbp<="011";
	end if;
	if (cc=180 and ll=198) then grbp<="011";
	end if;
	if (cc=236 and ll=198) then grbp<="011";
	end if;
	if (cc=72 and ll=199) then grbp<="011";
	end if;
	if (ll=199 and cc>=72 and cc<75) then grbp<="011";
	end if;
	if (cc=113 and ll=199) then grbp<="011";
	end if;
	if (cc=240 and ll=199) then grbp<="011";
	end if;
	if (cc=72 and ll=200) then grbp<="011";
	end if;
	if (ll=200 and cc>=72 and cc<74) then grbp<="011";
	end if;
	if (cc=104 and ll=200) then grbp<="011";
	end if;
	if (cc=107 and ll=200) then grbp<="011";
	end if;
	if (cc=239 and ll=200) then grbp<="011";
	end if;
	if (cc=71 and ll=201) then grbp<="011";
	end if;
	if (ll=201 and cc>=71 and cc<74) then grbp<="011";
	end if;
	if (cc=112 and ll=201) then grbp<="011";
	end if;
	if (cc=135 and ll=201) then grbp<="011";
	end if;
	if (cc=245 and ll=201) then grbp<="011";
	end if;
	if (cc=71 and ll=202) then grbp<="011";
	end if;
	if (ll=202 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (cc=104 and ll=202) then grbp<="011";
	end if;
	if (cc=236 and ll=202) then grbp<="011";
	end if;
	if (cc=70 and ll=203) then grbp<="011";
	end if;
	if (ll=203 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (cc=84 and ll=203) then grbp<="011";
	end if;
	if (ll=203 and cc>=84 and cc<86) then grbp<="011";
	end if;
	if (cc=114 and ll=203) then grbp<="011";
	end if;
	if (cc=138 and ll=203) then grbp<="011";
	end if;
	if (cc=240 and ll=203) then grbp<="011";
	end if;
	if (cc=244 and ll=203) then grbp<="011";
	end if;
	if (cc=70 and ll=204) then grbp<="011";
	end if;
	if (cc=84 and ll=204) then grbp<="011";
	end if;
	if (ll=204 and cc>=84 and cc<86) then grbp<="011";
	end if;
	if (ll=205 and cc>=84 and cc<86) then grbp<="011";
	end if;
	if (cc=79 and ll=206) then grbp<="011";
	end if;
	if (cc=85 and ll=206) then grbp<="011";
	end if;
	if (cc=239 and ll=206) then grbp<="011";
	end if;
	if (cc=69 and ll=207) then grbp<="011";
	end if;
	if (cc=79 and ll=207) then grbp<="011";
	end if;
	if (cc=85 and ll=207) then grbp<="011";
	end if;
	if (cc=101 and ll=207) then grbp<="011";
	end if;
	if (cc=112 and ll=207) then grbp<="011";
	end if;
	if (cc=241 and ll=207) then grbp<="011";
	end if;
	if (cc=69 and ll=208) then grbp<="011";
	end if;
	if (cc=83 and ll=208) then grbp<="011";
	end if;
	if (cc=85 and ll=208) then grbp<="011";
	end if;
	if (cc=243 and ll=208) then grbp<="011";
	end if;
	if (cc=69 and ll=209) then grbp<="011";
	end if;
	if (cc=78 and ll=209) then grbp<="011";
	end if;
	if (cc=82 and ll=209) then grbp<="011";
	end if;
	if (cc=85 and ll=209) then grbp<="011";
	end if;
	if (cc=103 and ll=209) then grbp<="011";
	end if;
	if (cc=243 and ll=209) then grbp<="011";
	end if;
	if (cc=69 and ll=210) then grbp<="011";
	end if;
	if (cc=78 and ll=210) then grbp<="011";
	end if;
	if (cc=82 and ll=210) then grbp<="011";
	end if;
	if (cc=85 and ll=210) then grbp<="011";
	end if;
	if (cc=134 and ll=210) then grbp<="011";
	end if;
	if (cc=77 and ll=211) then grbp<="011";
	end if;
	if (ll=211 and cc>=77 and cc<79) then grbp<="011";
	end if;
	if (cc=146 and ll=211) then grbp<="011";
	end if;
	if (cc=77 and ll=212) then grbp<="011";
	end if;
	if (cc=82 and ll=212) then grbp<="011";
	end if;
	if (cc=246 and ll=212) then grbp<="011";
	end if;
	if (cc=56 and ll=213) then grbp<="011";
	end if;
	if (cc=76 and ll=213) then grbp<="011";
	end if;
	if (ll=213 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=95 and ll=213) then grbp<="011";
	end if;
	if (cc=246 and ll=213) then grbp<="011";
	end if;
	if (cc=54 and ll=214) then grbp<="011";
	end if;
	if (ll=214 and cc>=54 and cc<56) then grbp<="011";
	end if;
	if (cc=95 and ll=214) then grbp<="011";
	end if;
	if (cc=245 and ll=214) then grbp<="011";
	end if;
	if (cc=73 and ll=215) then grbp<="011";
	end if;
	if (cc=76 and ll=215) then grbp<="011";
	end if;
	if (cc=81 and ll=215) then grbp<="011";
	end if;
	if (cc=96 and ll=215) then grbp<="011";
	end if;
	if (cc=53 and ll=216) then grbp<="011";
	end if;
	if (cc=72 and ll=216) then grbp<="011";
	end if;
	if (ll=216 and cc>=72 and cc<74) then grbp<="011";
	end if;
	if (cc=79 and ll=216) then grbp<="011";
	end if;
	if (cc=81 and ll=216) then grbp<="011";
	end if;
	if (cc=96 and ll=216) then grbp<="011";
	end if;
	if (ll=216 and cc>=96 and cc<98) then grbp<="011";
	end if;
	if (cc=243 and ll=216) then grbp<="011";
	end if;
	if (cc=72 and ll=217) then grbp<="011";
	end if;
	if (cc=75 and ll=217) then grbp<="011";
	end if;
	if (cc=79 and ll=217) then grbp<="011";
	end if;
	if (cc=81 and ll=217) then grbp<="011";
	end if;
	if (cc=97 and ll=217) then grbp<="011";
	end if;
	if (cc=134 and ll=217) then grbp<="011";
	end if;
	if (cc=181 and ll=217) then grbp<="011";
	end if;
	if (cc=71 and ll=218) then grbp<="011";
	end if;
	if (cc=79 and ll=218) then grbp<="011";
	end if;
	if (cc=97 and ll=218) then grbp<="011";
	end if;
	if (cc=135 and ll=218) then grbp<="011";
	end if;
	if (cc=240 and ll=218) then grbp<="011";
	end if;
	if (cc=74 and ll=219) then grbp<="011";
	end if;
	if (cc=78 and ll=219) then grbp<="011";
	end if;
	if (ll=219 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=163 and ll=219) then grbp<="011";
	end if;
	if (cc=165 and ll=219) then grbp<="011";
	end if;
	if (cc=70 and ll=220) then grbp<="011";
	end if;
	if (cc=78 and ll=220) then grbp<="011";
	end if;
	if (ll=220 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=90 and ll=220) then grbp<="011";
	end if;
	if (cc=163 and ll=220) then grbp<="011";
	end if;
	if (cc=181 and ll=220) then grbp<="011";
	end if;
	if (cc=238 and ll=220) then grbp<="011";
	end if;
	if (cc=78 and ll=221) then grbp<="011";
	end if;
	if (cc=81 and ll=221) then grbp<="011";
	end if;
	if (cc=90 and ll=221) then grbp<="011";
	end if;
	if (cc=164 and ll=221) then grbp<="011";
	end if;
	if (cc=240 and ll=221) then grbp<="011";
	end if;
	if (cc=68 and ll=222) then grbp<="011";
	end if;
	if (cc=78 and ll=222) then grbp<="011";
	end if;
	if (cc=81 and ll=222) then grbp<="011";
	end if;
	if (cc=90 and ll=222) then grbp<="011";
	end if;
	if (cc=240 and ll=222) then grbp<="011";
	end if;
	if (cc=249 and ll=222) then grbp<="011";
	end if;
	if (cc=68 and ll=223) then grbp<="011";
	end if;
	if (cc=78 and ll=223) then grbp<="011";
	end if;
	if (ll=223 and cc>=78 and cc<82) then grbp<="011";
	end if;
	if (cc=55 and ll=224) then grbp<="011";
	end if;
	if (cc=78 and ll=224) then grbp<="011";
	end if;
	if (ll=224 and cc>=78 and cc<82) then grbp<="011";
	end if;
	if (cc=54 and ll=225) then grbp<="011";
	end if;
	if (cc=78 and ll=225) then grbp<="011";
	end if;
	if (cc=81 and ll=225) then grbp<="011";
	end if;
	if (cc=131 and ll=225) then grbp<="011";
	end if;
	if (cc=158 and ll=225) then grbp<="011";
	end if;
	if (cc=239 and ll=225) then grbp<="011";
	end if;
	if (cc=54 and ll=226) then grbp<="011";
	end if;
	if (cc=78 and ll=226) then grbp<="011";
	end if;
	if (cc=81 and ll=226) then grbp<="011";
	end if;
	if (cc=128 and ll=226) then grbp<="011";
	end if;
	if (cc=130 and ll=226) then grbp<="011";
	end if;
	if (cc=158 and ll=226) then grbp<="011";
	end if;
	if (cc=162 and ll=226) then grbp<="011";
	end if;
	if (cc=51 and ll=227) then grbp<="011";
	end if;
	if (ll=227 and cc>=51 and cc<53) then grbp<="011";
	end if;
	if (ll=227 and cc>=66 and cc<68) then grbp<="011";
	end if;
	if (cc=80 and ll=227) then grbp<="011";
	end if;
	if (ll=227 and cc>=80 and cc<82) then grbp<="011";
	end if;
	if (ll=227 and cc>=129 and cc<131) then grbp<="011";
	end if;
	if (cc=159 and ll=227) then grbp<="011";
	end if;
	if (ll=227 and cc>=159 and cc<162) then grbp<="011";
	end if;
	if (cc=52 and ll=228) then grbp<="011";
	end if;
	if (cc=61 and ll=228) then grbp<="011";
	end if;
	if (cc=65 and ll=228) then grbp<="011";
	end if;
	if (ll=228 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=80 and ll=228) then grbp<="011";
	end if;
	if (ll=228 and cc>=80 and cc<83) then grbp<="011";
	end if;
	if (cc=138 and ll=228) then grbp<="011";
	end if;
	if (ll=228 and cc>=138 and cc<140) then grbp<="011";
	end if;
	if (cc=159 and ll=228) then grbp<="011";
	end if;
	if (ll=228 and cc>=159 and cc<162) then grbp<="011";
	end if;
	if (cc=51 and ll=229) then grbp<="011";
	end if;
	if (cc=61 and ll=229) then grbp<="011";
	end if;
	if (cc=63 and ll=229) then grbp<="011";
	end if;
	if (ll=229 and cc>=63 and cc<66) then grbp<="011";
	end if;
	if (ll=229 and cc>=78 and cc<83) then grbp<="011";
	end if;
	if (cc=51 and ll=230) then grbp<="011";
	end if;
	if (ll=230 and cc>=51 and cc<54) then grbp<="011";
	end if;
	if (ll=230 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=77 and ll=230) then grbp<="011";
	end if;
	if (ll=230 and cc>=77 and cc<83) then grbp<="011";
	end if;
	if (cc=50 and ll=231) then grbp<="011";
	end if;
	if (ll=231 and cc>=50 and cc<54) then grbp<="011";
	end if;
	if (cc=66 and ll=231) then grbp<="011";
	end if;
	if (cc=74 and ll=231) then grbp<="011";
	end if;
	if (cc=78 and ll=231) then grbp<="011";
	end if;
	if (ll=231 and cc>=78 and cc<84) then grbp<="011";
	end if;
	if (cc=136 and ll=231) then grbp<="011";
	end if;
	if (cc=182 and ll=231) then grbp<="011";
	end if;
	if (cc=49 and ll=232) then grbp<="011";
	end if;
	if (ll=232 and cc>=49 and cc<52) then grbp<="011";
	end if;
	if (ll=232 and cc>=62 and cc<64) then grbp<="011";
	end if;
	if (cc=77 and ll=232) then grbp<="011";
	end if;
	if (ll=232 and cc>=77 and cc<84) then grbp<="011";
	end if;
	if (cc=136 and ll=232) then grbp<="011";
	end if;
	if (ll=232 and cc>=136 and cc<139) then grbp<="011";
	end if;
	if (cc=182 and ll=232) then grbp<="011";
	end if;
	if (cc=46 and ll=233) then grbp<="011";
	end if;
	if (ll=233 and cc>=46 and cc<50) then grbp<="011";
	end if;
	if (ll=233 and cc>=64 and cc<69) then grbp<="011";
	end if;
	if (cc=77 and ll=233) then grbp<="011";
	end if;
	if (cc=79 and ll=233) then grbp<="011";
	end if;
	if (ll=233 and cc>=79 and cc<83) then grbp<="011";
	end if;
	if (cc=138 and ll=233) then grbp<="011";
	end if;
	if (ll=233 and cc>=138 and cc<141) then grbp<="011";
	end if;
	if (cc=180 and ll=233) then grbp<="011";
	end if;
	if (cc=45 and ll=234) then grbp<="011";
	end if;
	if (cc=64 and ll=234) then grbp<="011";
	end if;
	if (cc=66 and ll=234) then grbp<="011";
	end if;
	if (ll=234 and cc>=66 and cc<69) then grbp<="011";
	end if;
	if (cc=79 and ll=234) then grbp<="011";
	end if;
	if (ll=234 and cc>=79 and cc<84) then grbp<="011";
	end if;
	if (cc=133 and ll=234) then grbp<="011";
	end if;
	if (ll=234 and cc>=133 and cc<136) then grbp<="011";
	end if;
	if (cc=46 and ll=235) then grbp<="011";
	end if;
	if (cc=48 and ll=235) then grbp<="011";
	end if;
	if (cc=64 and ll=235) then grbp<="011";
	end if;
	if (ll=235 and cc>=64 and cc<68) then grbp<="011";
	end if;
	if (ll=235 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (cc=118 and ll=235) then grbp<="011";
	end if;
	if (cc=182 and ll=235) then grbp<="011";
	end if;
	if (cc=47 and ll=236) then grbp<="011";
	end if;
	if (cc=63 and ll=236) then grbp<="011";
	end if;
	if (cc=76 and ll=236) then grbp<="011";
	end if;
	if (ll=236 and cc>=76 and cc<80) then grbp<="011";
	end if;
	if (cc=83 and ll=236) then grbp<="011";
	end if;
	if (cc=126 and ll=236) then grbp<="011";
	end if;
	if (ll=236 and cc>=126 and cc<130) then grbp<="011";
	end if;
	if (cc=182 and ll=236) then grbp<="011";
	end if;
	if (cc=235 and ll=236) then grbp<="011";
	end if;
	if (cc=61 and ll=237) then grbp<="011";
	end if;
	if (ll=237 and cc>=61 and cc<64) then grbp<="011";
	end if;
	if (ll=237 and cc>=76 and cc<80) then grbp<="011";
	end if;
	if (cc=120 and ll=237) then grbp<="011";
	end if;
	if (cc=158 and ll=237) then grbp<="011";
	end if;
	if (cc=51 and ll=238) then grbp<="011";
	end if;
	if (ll=238 and cc>=51 and cc<53) then grbp<="011";
	end if;
	if (ll=238 and cc>=61 and cc<64) then grbp<="011";
	end if;
	if (cc=73 and ll=238) then grbp<="011";
	end if;
	if (cc=78 and ll=238) then grbp<="011";
	end if;
	if (cc=47 and ll=239) then grbp<="011";
	end if;
	if (ll=239 and cc>=47 and cc<51) then grbp<="011";
	end if;
	if (ll=239 and cc>=52 and cc<54) then grbp<="011";
	end if;
	if (cc=61 and ll=239) then grbp<="011";
	end if;
	if (cc=63 and ll=239) then grbp<="011";
	end if;
	if (cc=66 and ll=239) then grbp<="011";
	end if;
	if (cc=73 and ll=239) then grbp<="011";
	end if;
	if (cc=78 and ll=239) then grbp<="011";
	end if;
	if (ll=239 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=120 and ll=239) then grbp<="011";
	end if;
	if (cc=159 and ll=239) then grbp<="011";
	end if;
	if (cc=180 and ll=239) then grbp<="011";
	end if;
	if (cc=45 and ll=240) then grbp<="011";
	end if;
	if (ll=240 and cc>=45 and cc<48) then grbp<="011";
	end if;
	if (cc=59 and ll=240) then grbp<="011";
	end if;
	if (cc=61 and ll=240) then grbp<="011";
	end if;
	if (ll=240 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=73 and ll=240) then grbp<="011";
	end if;
	if (ll=240 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=240 and cc>=78 and cc<81) then grbp<="011";
	end if;
	if (cc=119 and ll=240) then grbp<="011";
	end if;
	if (cc=159 and ll=240) then grbp<="011";
	end if;
	if (cc=180 and ll=240) then grbp<="011";
	end if;
	if (cc=42 and ll=241) then grbp<="011";
	end if;
	if (ll=241 and cc>=42 and cc<46) then grbp<="011";
	end if;
	if (ll=241 and cc>=49 and cc<51) then grbp<="011";
	end if;
	if (ll=241 and cc>=61 and cc<66) then grbp<="011";
	end if;
	if (ll=241 and cc>=74 and cc<78) then grbp<="011";
	end if;
	if (cc=81 and ll=241) then grbp<="011";
	end if;
	if (cc=150 and ll=241) then grbp<="011";
	end if;
	if (cc=180 and ll=241) then grbp<="011";
	end if;
	if (cc=232 and ll=241) then grbp<="011";
	end if;
	if (cc=41 and ll=242) then grbp<="011";
	end if;
	if (cc=58 and ll=242) then grbp<="011";
	end if;
	if (cc=61 and ll=242) then grbp<="011";
	end if;
	if (cc=63 and ll=242) then grbp<="011";
	end if;
	if (ll=242 and cc>=63 and cc<66) then grbp<="011";
	end if;
	if (ll=242 and cc>=76 and cc<80) then grbp<="011";
	end if;
	if (cc=180 and ll=242) then grbp<="011";
	end if;
	if (cc=183 and ll=242) then grbp<="011";
	end if;
	if (cc=40 and ll=243) then grbp<="011";
	end if;
	if (cc=43 and ll=243) then grbp<="011";
	end if;
	if (ll=243 and cc>=43 and cc<46) then grbp<="011";
	end if;
	if (cc=62 and ll=243) then grbp<="011";
	end if;
	if (ll=243 and cc>=62 and cc<65) then grbp<="011";
	end if;
	if (ll=243 and cc>=77 and cc<79) then grbp<="011";
	end if;
	if (cc=139 and ll=243) then grbp<="011";
	end if;
	if (cc=39 and ll=244) then grbp<="011";
	end if;
	if (cc=43 and ll=244) then grbp<="011";
	end if;
	if (ll=244 and cc>=43 and cc<46) then grbp<="011";
	end if;
	if (ll=244 and cc>=60 and cc<65) then grbp<="011";
	end if;
	if (cc=150 and ll=244) then grbp<="011";
	end if;
	if (cc=43 and ll=245) then grbp<="011";
	end if;
	if (cc=45 and ll=245) then grbp<="011";
	end if;
	if (ll=245 and cc>=45 and cc<47) then grbp<="011";
	end if;
	if (cc=60 and ll=245) then grbp<="011";
	end if;
	if (ll=245 and cc>=60 and cc<65) then grbp<="011";
	end if;
	if (ll=246 and cc>=56 and cc<58) then grbp<="011";
	end if;
	if (ll=246 and cc>=60 and cc<63) then grbp<="011";
	end if;
	if (cc=49 and ll=247) then grbp<="011";
	end if;
	if (cc=56 and ll=247) then grbp<="011";
	end if;
	if (cc=60 and ll=247) then grbp<="011";
	end if;
	if (cc=62 and ll=247) then grbp<="011";
	end if;
	if (cc=48 and ll=248) then grbp<="011";
	end if;
	if (ll=248 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (cc=59 and ll=248) then grbp<="011";
	end if;
	if (cc=62 and ll=248) then grbp<="011";
	end if;
	if (cc=160 and ll=248) then grbp<="011";
	end if;
	if (cc=214 and ll=248) then grbp<="011";
	end if;
	if (cc=46 and ll=249) then grbp<="011";
	end if;
	if (ll=249 and cc>=46 and cc<49) then grbp<="011";
	end if;
	if (ll=249 and cc>=54 and cc<56) then grbp<="011";
	end if;
	if (ll=249 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=182 and ll=249) then grbp<="011";
	end if;
	if (cc=45 and ll=250) then grbp<="011";
	end if;
	if (ll=250 and cc>=45 and cc<48) then grbp<="011";
	end if;
	if (cc=60 and ll=250) then grbp<="011";
	end if;
	if (ll=250 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (cc=44 and ll=251) then grbp<="011";
	end if;
	if (cc=46 and ll=251) then grbp<="011";
	end if;
	if (cc=50 and ll=251) then grbp<="011";
	end if;
	if (cc=53 and ll=251) then grbp<="011";
	end if;
	if (cc=61 and ll=251) then grbp<="011";
	end if;
	if (cc=162 and ll=251) then grbp<="011";
	end if;
	if (cc=184 and ll=251) then grbp<="011";
	end if;
	if (cc=36 and ll=252) then grbp<="011";
	end if;
	if (cc=43 and ll=252) then grbp<="011";
	end if;
	if (ll=252 and cc>=43 and cc<45) then grbp<="011";
	end if;
	if (ll=252 and cc>=49 and cc<51) then grbp<="011";
	end if;
	if (ll=252 and cc>=52 and cc<54) then grbp<="011";
	end if;
	if (cc=63 and ll=252) then grbp<="011";
	end if;
	if (cc=151 and ll=252) then grbp<="011";
	end if;
	if (cc=183 and ll=252) then grbp<="011";
	end if;
	if (ll=252 and cc>=183 and cc<185) then grbp<="011";
	end if;
	if (cc=41 and ll=253) then grbp<="011";
	end if;
	if (ll=253 and cc>=41 and cc<43) then grbp<="011";
	end if;
	if (cc=49 and ll=253) then grbp<="011";
	end if;
	if (ll=253 and cc>=49 and cc<51) then grbp<="011";
	end if;
	if (cc=56 and ll=253) then grbp<="011";
	end if;
	if (cc=60 and ll=253) then grbp<="011";
	end if;
	if (ll=253 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (cc=83 and ll=253) then grbp<="011";
	end if;
	if (cc=183 and ll=253) then grbp<="011";
	end if;
	if (cc=36 and ll=254) then grbp<="011";
	end if;
	if (cc=40 and ll=254) then grbp<="011";
	end if;
	if (cc=43 and ll=254) then grbp<="011";
	end if;
	if (cc=48 and ll=254) then grbp<="011";
	end if;
	if (cc=51 and ll=254) then grbp<="011";
	end if;
	if (cc=56 and ll=254) then grbp<="011";
	end if;
	if (cc=60 and ll=254) then grbp<="011";
	end if;
	if (ll=254 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (ll=254 and cc>=183 and cc<185) then grbp<="011";
	end if;
	if (cc=39 and ll=255) then grbp<="011";
	end if;
	if (cc=41 and ll=255) then grbp<="011";
	end if;
	if (cc=43 and ll=255) then grbp<="011";
	end if;
	if (cc=48 and ll=255) then grbp<="011";
	end if;
	if (ll=255 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (cc=56 and ll=255) then grbp<="011";
	end if;
	if (cc=60 and ll=255) then grbp<="011";
	end if;
	if (ll=255 and cc>=60 and cc<64) then grbp<="011";
	end if;
	if (cc=183 and ll=255) then grbp<="011";
	end if;
	if (cc=37 and ll=256) then grbp<="011";
	end if;
	if (cc=40 and ll=256) then grbp<="011";
	end if;
	if (cc=42 and ll=256) then grbp<="011";
	end if;
	if (ll=256 and cc>=42 and cc<44) then grbp<="011";
	end if;
	if (ll=256 and cc>=47 and cc<49) then grbp<="011";
	end if;
	if (cc=57 and ll=256) then grbp<="011";
	end if;
	if (cc=59 and ll=256) then grbp<="011";
	end if;
	if (ll=256 and cc>=59 and cc<63) then grbp<="011";
	end if;
	if (cc=82 and ll=256) then grbp<="011";
	end if;
	if (cc=151 and ll=256) then grbp<="011";
	end if;
	if (cc=38 and ll=257) then grbp<="011";
	end if;
	if (ll=257 and cc>=38 and cc<40) then grbp<="011";
	end if;
	if (cc=47 and ll=257) then grbp<="011";
	end if;
	if (ll=257 and cc>=47 and cc<49) then grbp<="011";
	end if;
	if (cc=57 and ll=257) then grbp<="011";
	end if;
	if (cc=59 and ll=257) then grbp<="011";
	end if;
	if (ll=257 and cc>=59 and cc<63) then grbp<="011";
	end if;
	if (cc=151 and ll=257) then grbp<="011";
	end if;
	if (cc=159 and ll=257) then grbp<="011";
	end if;
	if (cc=181 and ll=257) then grbp<="011";
	end if;
	if (cc=38 and ll=258) then grbp<="011";
	end if;
	if (ll=258 and cc>=38 and cc<40) then grbp<="011";
	end if;
	if (cc=55 and ll=258) then grbp<="011";
	end if;
	if (cc=57 and ll=258) then grbp<="011";
	end if;
	if (cc=59 and ll=258) then grbp<="011";
	end if;
	if (ll=258 and cc>=59 and cc<62) then grbp<="011";
	end if;
	if (cc=181 and ll=258) then grbp<="011";
	end if;
	if (cc=39 and ll=259) then grbp<="011";
	end if;
	if (ll=259 and cc>=39 and cc<44) then grbp<="011";
	end if;
	if (cc=56 and ll=259) then grbp<="011";
	end if;
	if (ll=259 and cc>=56 and cc<58) then grbp<="011";
	end if;
	if (cc=61 and ll=259) then grbp<="011";
	end if;
	if (cc=64 and ll=259) then grbp<="011";
	end if;
	if (cc=80 and ll=259) then grbp<="011";
	end if;
	if (cc=39 and ll=260) then grbp<="011";
	end if;
	if (cc=41 and ll=260) then grbp<="011";
	end if;
	if (ll=260 and cc>=41 and cc<44) then grbp<="011";
	end if;
	if (cc=56 and ll=260) then grbp<="011";
	end if;
	if (cc=59 and ll=260) then grbp<="011";
	end if;
	if (cc=61 and ll=260) then grbp<="011";
	end if;
	if (cc=49 and ll=261) then grbp<="011";
	end if;
	if (cc=56 and ll=261) then grbp<="011";
	end if;
	if (cc=59 and ll=261) then grbp<="011";
	end if;
	if (cc=61 and ll=261) then grbp<="011";
	end if;
	if (cc=128 and ll=261) then grbp<="011";
	end if;
	if (cc=183 and ll=261) then grbp<="011";
	end if;
	if (cc=37 and ll=262) then grbp<="011";
	end if;
	if (ll=262 and cc>=37 and cc<39) then grbp<="011";
	end if;
	if (cc=55 and ll=262) then grbp<="011";
	end if;
	if (ll=262 and cc>=55 and cc<57) then grbp<="011";
	end if;
	if (cc=61 and ll=262) then grbp<="011";
	end if;
	if (cc=98 and ll=262) then grbp<="011";
	end if;
	if (cc=36 and ll=263) then grbp<="011";
	end if;
	if (ll=263 and cc>=36 and cc<38) then grbp<="011";
	end if;
	if (ll=263 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (cc=59 and ll=263) then grbp<="011";
	end if;
	if (cc=61 and ll=263) then grbp<="011";
	end if;
	if (cc=65 and ll=263) then grbp<="011";
	end if;
	if (cc=90 and ll=263) then grbp<="011";
	end if;
	if (cc=128 and ll=263) then grbp<="011";
	end if;
	if (cc=36 and ll=264) then grbp<="011";
	end if;
	if (cc=48 and ll=264) then grbp<="011";
	end if;
	if (ll=264 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (cc=59 and ll=264) then grbp<="011";
	end if;
	if (cc=61 and ll=264) then grbp<="011";
	end if;
	if (cc=65 and ll=264) then grbp<="011";
	end if;
	if (cc=95 and ll=264) then grbp<="011";
	end if;
	if (cc=134 and ll=264) then grbp<="011";
	end if;
	if (cc=35 and ll=265) then grbp<="011";
	end if;
	if (cc=47 and ll=265) then grbp<="011";
	end if;
	if (ll=265 and cc>=47 and cc<49) then grbp<="011";
	end if;
	if (cc=59 and ll=265) then grbp<="011";
	end if;
	if (cc=63 and ll=265) then grbp<="011";
	end if;
	if (cc=81 and ll=265) then grbp<="011";
	end if;
	if (cc=47 and ll=266) then grbp<="011";
	end if;
	if (ll=266 and cc>=47 and cc<50) then grbp<="011";
	end if;
	if (ll=266 and cc>=54 and cc<56) then grbp<="011";
	end if;
	if (cc=63 and ll=266) then grbp<="011";
	end if;
	if (cc=65 and ll=266) then grbp<="011";
	end if;
	if (cc=130 and ll=266) then grbp<="011";
	end if;
	if (cc=42 and ll=267) then grbp<="011";
	end if;
	if (cc=47 and ll=267) then grbp<="011";
	end if;
	if (ll=267 and cc>=47 and cc<50) then grbp<="011";
	end if;
	if (cc=59 and ll=267) then grbp<="011";
	end if;
	if (cc=65 and ll=267) then grbp<="011";
	end if;
	if (cc=80 and ll=267) then grbp<="011";
	end if;
	if (cc=46 and ll=268) then grbp<="011";
	end if;
	if (cc=48 and ll=268) then grbp<="011";
	end if;
	if (ll=268 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (ll=268 and cc>=59 and cc<61) then grbp<="011";
	end if;
	if (cc=182 and ll=268) then grbp<="011";
	end if;
	if (cc=185 and ll=268) then grbp<="011";
	end if;
	if (cc=48 and ll=269) then grbp<="011";
	end if;
	if (cc=54 and ll=269) then grbp<="011";
	end if;
	if (cc=59 and ll=269) then grbp<="011";
	end if;
	if (cc=62 and ll=269) then grbp<="011";
	end if;
	if (cc=66 and ll=269) then grbp<="011";
	end if;
	if (cc=134 and ll=269) then grbp<="011";
	end if;
	if (cc=53 and ll=270) then grbp<="011";
	end if;
	if (ll=270 and cc>=53 and cc<55) then grbp<="011";
	end if;
	if (cc=62 and ll=270) then grbp<="011";
	end if;
	if (cc=66 and ll=270) then grbp<="011";
	end if;
	if (cc=79 and ll=270) then grbp<="011";
	end if;
	if (cc=53 and ll=271) then grbp<="011";
	end if;
	if (ll=271 and cc>=53 and cc<55) then grbp<="011";
	end if;
	if (ll=271 and cc>=59 and cc<61) then grbp<="011";
	end if;
	if (cc=64 and ll=271) then grbp<="011";
	end if;
	if (cc=79 and ll=271) then grbp<="011";
	end if;
	if (cc=184 and ll=271) then grbp<="011";
	end if;
	if (cc=52 and ll=272) then grbp<="011";
	end if;
	if (ll=272 and cc>=52 and cc<54) then grbp<="011";
	end if;
	if (ll=272 and cc>=59 and cc<61) then grbp<="011";
	end if;
	if (ll=272 and cc>=62 and cc<65) then grbp<="011";
	end if;
	if (cc=151 and ll=272) then grbp<="011";
	end if;
	if (cc=184 and ll=272) then grbp<="011";
	end if;
	if (cc=52 and ll=273) then grbp<="011";
	end if;
	if (cc=60 and ll=273) then grbp<="011";
	end if;
	if (cc=62 and ll=273) then grbp<="011";
	end if;
	if (cc=65 and ll=273) then grbp<="011";
	end if;
	if (ll=273 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=150 and ll=273) then grbp<="011";
	end if;
	if (cc=184 and ll=273) then grbp<="011";
	end if;
	if (cc=213 and ll=273) then grbp<="011";
	end if;
	if (cc=51 and ll=274) then grbp<="011";
	end if;
	if (cc=59 and ll=274) then grbp<="011";
	end if;
	if (ll=274 and cc>=59 and cc<61) then grbp<="011";
	end if;
	if (cc=65 and ll=274) then grbp<="011";
	end if;
	if (ll=274 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=184 and ll=274) then grbp<="011";
	end if;
	if (cc=42 and ll=275) then grbp<="011";
	end if;
	if (cc=51 and ll=275) then grbp<="011";
	end if;
	if (cc=59 and ll=275) then grbp<="011";
	end if;
	if (ll=275 and cc>=59 and cc<63) then grbp<="011";
	end if;
	if (cc=67 and ll=275) then grbp<="011";
	end if;
	if (cc=84 and ll=275) then grbp<="011";
	end if;
	if (cc=42 and ll=276) then grbp<="011";
	end if;
	if (cc=50 and ll=276) then grbp<="011";
	end if;
	if (cc=59 and ll=276) then grbp<="011";
	end if;
	if (ll=276 and cc>=59 and cc<63) then grbp<="011";
	end if;
	if (cc=67 and ll=276) then grbp<="011";
	end if;
	if (cc=41 and ll=277) then grbp<="011";
	end if;
	if (ll=277 and cc>=41 and cc<43) then grbp<="011";
	end if;
	if (ll=277 and cc>=49 and cc<51) then grbp<="011";
	end if;
	if (cc=61 and ll=277) then grbp<="011";
	end if;
	if (ll=277 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=277 and cc>=65 and cc<68) then grbp<="011";
	end if;
	if (cc=40 and ll=278) then grbp<="011";
	end if;
	if (ll=278 and cc>=40 and cc<42) then grbp<="011";
	end if;
	if (ll=278 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (ll=278 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=278 and cc>=64 and cc<68) then grbp<="011";
	end if;
	if (ll=278 and cc>=80 and cc<83) then grbp<="011";
	end if;
	if (cc=48 and ll=279) then grbp<="011";
	end if;
	if (ll=279 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (ll=279 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=279 and cc>=65 and cc<69) then grbp<="011";
	end if;
	if (cc=183 and ll=279) then grbp<="011";
	end if;
	if (cc=40 and ll=280) then grbp<="011";
	end if;
	if (cc=42 and ll=280) then grbp<="011";
	end if;
	if (cc=47 and ll=280) then grbp<="011";
	end if;
	if (ll=280 and cc>=47 and cc<49) then grbp<="011";
	end if;
	if (ll=280 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=280 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=79 and ll=280) then grbp<="011";
	end if;
	if (cc=81 and ll=280) then grbp<="011";
	end if;
	if (cc=39 and ll=281) then grbp<="011";
	end if;
	if (cc=47 and ll=281) then grbp<="011";
	end if;
	if (ll=281 and cc>=47 and cc<49) then grbp<="011";
	end if;
	if (cc=65 and ll=281) then grbp<="011";
	end if;
	if (ll=281 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=39 and ll=282) then grbp<="011";
	end if;
	if (cc=46 and ll=282) then grbp<="011";
	end if;
	if (ll=282 and cc>=46 and cc<48) then grbp<="011";
	end if;
	if (cc=65 and ll=282) then grbp<="011";
	end if;
	if (ll=282 and cc>=65 and cc<69) then grbp<="011";
	end if;
	if (cc=38 and ll=283) then grbp<="011";
	end if;
	if (cc=46 and ll=283) then grbp<="011";
	end if;
	if (ll=283 and cc>=46 and cc<48) then grbp<="011";
	end if;
	if (cc=65 and ll=283) then grbp<="011";
	end if;
	if (ll=283 and cc>=65 and cc<71) then grbp<="011";
	end if;
	if (cc=38 and ll=284) then grbp<="011";
	end if;
	if (cc=42 and ll=284) then grbp<="011";
	end if;
	if (cc=47 and ll=284) then grbp<="011";
	end if;
	if (cc=66 and ll=284) then grbp<="011";
	end if;
	if (ll=284 and cc>=66 and cc<70) then grbp<="011";
	end if;
	if (cc=37 and ll=285) then grbp<="011";
	end if;
	if (cc=63 and ll=285) then grbp<="011";
	end if;
	if (cc=66 and ll=285) then grbp<="011";
	end if;
	if (cc=68 and ll=285) then grbp<="011";
	end if;
	if (cc=70 and ll=285) then grbp<="011";
	end if;
	if (cc=76 and ll=285) then grbp<="011";
	end if;
	if (ll=285 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=143 and ll=285) then grbp<="011";
	end if;
	if (cc=37 and ll=286) then grbp<="011";
	end if;
	if (cc=46 and ll=286) then grbp<="011";
	end if;
	if (cc=56 and ll=286) then grbp<="011";
	end if;
	if (cc=67 and ll=286) then grbp<="011";
	end if;
	if (ll=286 and cc>=67 and cc<69) then grbp<="011";
	end if;
	if (cc=46 and ll=287) then grbp<="011";
	end if;
	if (ll=287 and cc>=46 and cc<48) then grbp<="011";
	end if;
	if (cc=69 and ll=287) then grbp<="011";
	end if;
	if (ll=287 and cc>=69 and cc<71) then grbp<="011";
	end if;
	if (cc=151 and ll=287) then grbp<="011";
	end if;
	if (ll=287 and cc>=151 and cc<153) then grbp<="011";
	end if;
	if (cc=41 and ll=288) then grbp<="011";
	end if;
	if (cc=47 and ll=288) then grbp<="011";
	end if;
	if (cc=57 and ll=288) then grbp<="011";
	end if;
	if (cc=59 and ll=288) then grbp<="011";
	end if;
	if (cc=64 and ll=288) then grbp<="011";
	end if;
	if (cc=69 and ll=288) then grbp<="011";
	end if;
	if (ll=288 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=57 and ll=289) then grbp<="011";
	end if;
	if (cc=60 and ll=289) then grbp<="011";
	end if;
	if (cc=65 and ll=289) then grbp<="011";
	end if;
	if (cc=69 and ll=289) then grbp<="011";
	end if;
	if (ll=289 and cc>=69 and cc<76) then grbp<="011";
	end if;
	if (cc=35 and ll=290) then grbp<="011";
	end if;
	if (cc=40 and ll=290) then grbp<="011";
	end if;
	if (cc=57 and ll=290) then grbp<="011";
	end if;
	if (ll=290 and cc>=57 and cc<61) then grbp<="011";
	end if;
	if (ll=290 and cc>=65 and cc<68) then grbp<="011";
	end if;
	if (cc=72 and ll=290) then grbp<="011";
	end if;
	if (cc=75 and ll=290) then grbp<="011";
	end if;
	if (cc=85 and ll=290) then grbp<="011";
	end if;
	if (cc=185 and ll=290) then grbp<="011";
	end if;
	if (ll=290 and cc>=185 and cc<187) then grbp<="011";
	end if;
	if (cc=40 and ll=291) then grbp<="011";
	end if;
	if (ll=291 and cc>=40 and cc<42) then grbp<="011";
	end if;
	if (ll=291 and cc>=57 and cc<62) then grbp<="011";
	end if;
	if (ll=291 and cc>=66 and cc<68) then grbp<="011";
	end if;
	if (cc=185 and ll=291) then grbp<="011";
	end if;
	if (cc=34 and ll=292) then grbp<="011";
	end if;
	if (cc=39 and ll=292) then grbp<="011";
	end if;
	if (ll=292 and cc>=39 and cc<42) then grbp<="011";
	end if;
	if (ll=292 and cc>=56 and cc<64) then grbp<="011";
	end if;
	if (cc=185 and ll=292) then grbp<="011";
	end if;
	if (cc=34 and ll=293) then grbp<="011";
	end if;
	if (cc=39 and ll=293) then grbp<="011";
	end if;
	if (ll=293 and cc>=39 and cc<41) then grbp<="011";
	end if;
	if (ll=293 and cc>=56 and cc<65) then grbp<="011";
	end if;
	if (ll=293 and cc>=66 and cc<68) then grbp<="011";
	end if;
	if (ll=293 and cc>=148 and cc<152) then grbp<="011";
	end if;
	if (cc=39 and ll=294) then grbp<="011";
	end if;
	if (cc=56 and ll=294) then grbp<="011";
	end if;
	if (cc=58 and ll=294) then grbp<="011";
	end if;
	if (cc=64 and ll=294) then grbp<="011";
	end if;
	if (cc=68 and ll=294) then grbp<="011";
	end if;
	if (cc=71 and ll=294) then grbp<="011";
	end if;
	if (ll=294 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (cc=143 and ll=294) then grbp<="011";
	end if;
	if (ll=294 and cc>=143 and cc<147) then grbp<="011";
	end if;
	if (cc=32 and ll=295) then grbp<="011";
	end if;
	if (ll=295 and cc>=32 and cc<34) then grbp<="011";
	end if;
	if (cc=56 and ll=295) then grbp<="011";
	end if;
	if (cc=58 and ll=295) then grbp<="011";
	end if;
	if (cc=61 and ll=295) then grbp<="011";
	end if;
	if (ll=295 and cc>=61 and cc<64) then grbp<="011";
	end if;
	if (ll=295 and cc>=70 and cc<73) then grbp<="011";
	end if;
	if (cc=151 and ll=295) then grbp<="011";
	end if;
	if (cc=184 and ll=295) then grbp<="011";
	end if;
	if (cc=32 and ll=296) then grbp<="011";
	end if;
	if (cc=38 and ll=296) then grbp<="011";
	end if;
	if (cc=45 and ll=296) then grbp<="011";
	end if;
	if (cc=54 and ll=296) then grbp<="011";
	end if;
	if (cc=56 and ll=296) then grbp<="011";
	end if;
	if (cc=58 and ll=296) then grbp<="011";
	end if;
	if (cc=62 and ll=296) then grbp<="011";
	end if;
	if (ll=296 and cc>=62 and cc<64) then grbp<="011";
	end if;
	if (ll=296 and cc>=69 and cc<73) then grbp<="011";
	end if;
	if (cc=30 and ll=297) then grbp<="011";
	end if;
	if (ll=297 and cc>=30 and cc<33) then grbp<="011";
	end if;
	if (cc=45 and ll=297) then grbp<="011";
	end if;
	if (cc=51 and ll=297) then grbp<="011";
	end if;
	if (cc=56 and ll=297) then grbp<="011";
	end if;
	if (cc=58 and ll=297) then grbp<="011";
	end if;
	if (cc=63 and ll=297) then grbp<="011";
	end if;
	if (ll=297 and cc>=63 and cc<65) then grbp<="011";
	end if;
	if (ll=297 and cc>=70 and cc<74) then grbp<="011";
	end if;
	if (cc=144 and ll=297) then grbp<="011";
	end if;
	if (cc=146 and ll=297) then grbp<="011";
	end if;
	if (ll=297 and cc>=146 and cc<149) then grbp<="011";
	end if;
	if (cc=37 and ll=298) then grbp<="011";
	end if;
	if (cc=51 and ll=298) then grbp<="011";
	end if;
	if (cc=58 and ll=298) then grbp<="011";
	end if;
	if (cc=64 and ll=298) then grbp<="011";
	end if;
	if (ll=298 and cc>=64 and cc<66) then grbp<="011";
	end if;
	if (ll=298 and cc>=70 and cc<74) then grbp<="011";
	end if;
	if (ll=298 and cc>=144 and cc<148) then grbp<="011";
	end if;
	if (ll=298 and cc>=149 and cc<151) then grbp<="011";
	end if;
	if (cc=45 and ll=299) then grbp<="011";
	end if;
	if (cc=51 and ll=299) then grbp<="011";
	end if;
	if (cc=57 and ll=299) then grbp<="011";
	end if;
	if (ll=299 and cc>=57 and cc<60) then grbp<="011";
	end if;
	if (ll=299 and cc>=64 and cc<67) then grbp<="011";
	end if;
	if (ll=299 and cc>=69 and cc<71) then grbp<="011";
	end if;
	if (ll=299 and cc>=72 and cc<74) then grbp<="011";
	end if;
	if (ll=299 and cc>=145 and cc<147) then grbp<="011";
	end if;
	if (cc=44 and ll=300) then grbp<="011";
	end if;
	if (ll=300 and cc>=44 and cc<46) then grbp<="011";
	end if;
	if (cc=57 and ll=300) then grbp<="011";
	end if;
	if (cc=59 and ll=300) then grbp<="011";
	end if;
	if (cc=62 and ll=300) then grbp<="011";
	end if;
	if (cc=65 and ll=300) then grbp<="011";
	end if;
	if (ll=300 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (ll=300 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (cc=36 and ll=301) then grbp<="011";
	end if;
	if (cc=44 and ll=301) then grbp<="011";
	end if;
	if (ll=301 and cc>=44 and cc<46) then grbp<="011";
	end if;
	if (cc=61 and ll=301) then grbp<="011";
	end if;
	if (ll=301 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=301 and cc>=66 and cc<72) then grbp<="011";
	end if;
	if (cc=44 and ll=302) then grbp<="011";
	end if;
	if (ll=302 and cc>=44 and cc<46) then grbp<="011";
	end if;
	if (cc=59 and ll=302) then grbp<="011";
	end if;
	if (ll=302 and cc>=59 and cc<63) then grbp<="011";
	end if;
	if (ll=302 and cc>=66 and cc<69) then grbp<="011";
	end if;
	if (cc=73 and ll=302) then grbp<="011";
	end if;
	if (ll=302 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (cc=55 and ll=303) then grbp<="011";
	end if;
	if (cc=57 and ll=303) then grbp<="011";
	end if;
	if (cc=60 and ll=303) then grbp<="011";
	end if;
	if (ll=303 and cc>=60 and cc<63) then grbp<="011";
	end if;
	if (cc=70 and ll=303) then grbp<="011";
	end if;
	if (cc=72 and ll=303) then grbp<="011";
	end if;
	if (cc=74 and ll=303) then grbp<="011";
	end if;
	if (ll=303 and cc>=74 and cc<76) then grbp<="011";
	end if;
	if (cc=44 and ll=304) then grbp<="011";
	end if;
	if (cc=55 and ll=304) then grbp<="011";
	end if;
	if (cc=61 and ll=304) then grbp<="011";
	end if;
	if (ll=304 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=304 and cc>=66 and cc<70) then grbp<="011";
	end if;
	if (cc=74 and ll=304) then grbp<="011";
	end if;
	if (ll=304 and cc>=74 and cc<76) then grbp<="011";
	end if;
	if (cc=58 and ll=305) then grbp<="011";
	end if;
	if (cc=61 and ll=305) then grbp<="011";
	end if;
	if (ll=305 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=305 and cc>=65 and cc<70) then grbp<="011";
	end if;
	if (cc=74 and ll=305) then grbp<="011";
	end if;
	if (cc=44 and ll=306) then grbp<="011";
	end if;
	if (cc=57 and ll=306) then grbp<="011";
	end if;
	if (ll=306 and cc>=57 and cc<59) then grbp<="011";
	end if;
	if (ll=306 and cc>=60 and cc<66) then grbp<="011";
	end if;
	if (ll=306 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (ll=306 and cc>=72 and cc<76) then grbp<="011";
	end if;
	if (cc=36 and ll=307) then grbp<="011";
	end if;
	if (cc=57 and ll=307) then grbp<="011";
	end if;
	if (ll=307 and cc>=57 and cc<60) then grbp<="011";
	end if;
	if (ll=307 and cc>=62 and cc<66) then grbp<="011";
	end if;
	if (ll=307 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (cc=74 and ll=307) then grbp<="011";
	end if;
	if (cc=36 and ll=308) then grbp<="011";
	end if;
	if (cc=55 and ll=308) then grbp<="011";
	end if;
	if (ll=308 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (cc=62 and ll=308) then grbp<="011";
	end if;
	if (ll=308 and cc>=62 and cc<65) then grbp<="011";
	end if;
	if (ll=308 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (cc=74 and ll=308) then grbp<="011";
	end if;
	if (cc=55 and ll=309) then grbp<="011";
	end if;
	if (ll=309 and cc>=55 and cc<61) then grbp<="011";
	end if;
	if (ll=309 and cc>=62 and cc<65) then grbp<="011";
	end if;
	if (ll=309 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (cc=74 and ll=309) then grbp<="011";
	end if;
	if (cc=55 and ll=310) then grbp<="011";
	end if;
	if (ll=310 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=310 and cc>=59 and cc<66) then grbp<="011";
	end if;
	if (cc=72 and ll=310) then grbp<="011";
	end if;
	if (cc=74 and ll=310) then grbp<="011";
	end if;
	if (cc=137 and ll=310) then grbp<="011";
	end if;
	if (cc=55 and ll=311) then grbp<="011";
	end if;
	if (ll=311 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=311 and cc>=59 and cc<67) then grbp<="011";
	end if;
	if (cc=72 and ll=311) then grbp<="011";
	end if;
	if (cc=75 and ll=311) then grbp<="011";
	end if;
	if (cc=77 and ll=311) then grbp<="011";
	end if;
	if (cc=136 and ll=311) then grbp<="011";
	end if;
	if (cc=139 and ll=311) then grbp<="011";
	end if;
	if (cc=149 and ll=311) then grbp<="011";
	end if;
	if (cc=55 and ll=312) then grbp<="011";
	end if;
	if (cc=57 and ll=312) then grbp<="011";
	end if;
	if (cc=61 and ll=312) then grbp<="011";
	end if;
	if (ll=312 and cc>=61 and cc<67) then grbp<="011";
	end if;
	if (cc=75 and ll=312) then grbp<="011";
	end if;
	if (cc=77 and ll=312) then grbp<="011";
	end if;
	if (cc=43 and ll=313) then grbp<="011";
	end if;
	if (cc=55 and ll=313) then grbp<="011";
	end if;
	if (cc=57 and ll=313) then grbp<="011";
	end if;
	if (cc=61 and ll=313) then grbp<="011";
	end if;
	if (ll=313 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=313 and cc>=64 and cc<68) then grbp<="011";
	end if;
	if (cc=72 and ll=313) then grbp<="011";
	end if;
	if (cc=135 and ll=313) then grbp<="011";
	end if;
	if (cc=149 and ll=313) then grbp<="011";
	end if;
	if (cc=43 and ll=314) then grbp<="011";
	end if;
	if (cc=55 and ll=314) then grbp<="011";
	end if;
	if (ll=314 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=314 and cc>=62 and cc<73) then grbp<="011";
	end if;
	if (cc=55 and ll=315) then grbp<="011";
	end if;
	if (ll=315 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=315 and cc>=63 and cc<73) then grbp<="011";
	end if;
	if (cc=55 and ll=316) then grbp<="011";
	end if;
	if (ll=316 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=316 and cc>=63 and cc<66) then grbp<="011";
	end if;
	if (ll=316 and cc>=67 and cc<73) then grbp<="011";
	end if;
	if (cc=55 and ll=317) then grbp<="011";
	end if;
	if (ll=317 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (ll=317 and cc>=63 and cc<67) then grbp<="011";
	end if;
	if (ll=317 and cc>=68 and cc<72) then grbp<="011";
	end if;
	if (cc=136 and ll=317) then grbp<="011";
	end if;
	if (cc=210 and ll=317) then grbp<="011";
	end if;
	if (cc=55 and ll=318) then grbp<="011";
	end if;
	if (ll=318 and cc>=55 and cc<58) then grbp<="011";
	end if;
	if (cc=65 and ll=318) then grbp<="011";
	end if;
	if (ll=318 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (ll=318 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=75 and ll=318) then grbp<="011";
	end if;
	if (cc=137 and ll=318) then grbp<="011";
	end if;
	if (cc=139 and ll=318) then grbp<="011";
	end if;
	if (cc=36 and ll=319) then grbp<="011";
	end if;
	if (cc=57 and ll=319) then grbp<="011";
	end if;
	if (cc=63 and ll=319) then grbp<="011";
	end if;
	if (ll=319 and cc>=63 and cc<66) then grbp<="011";
	end if;
	if (ll=319 and cc>=67 and cc<72) then grbp<="011";
	end if;
	if (ll=319 and cc>=73 and cc<77) then grbp<="011";
	end if;
	if (cc=58 and ll=320) then grbp<="011";
	end if;
	if (cc=64 and ll=320) then grbp<="011";
	end if;
	if (ll=320 and cc>=64 and cc<66) then grbp<="011";
	end if;
	if (ll=320 and cc>=67 and cc<71) then grbp<="011";
	end if;
	if (ll=320 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (cc=209 and ll=320) then grbp<="011";
	end if;
	if (cc=34 and ll=321) then grbp<="011";
	end if;
	if (cc=57 and ll=321) then grbp<="011";
	end if;
	if (ll=321 and cc>=57 and cc<61) then grbp<="011";
	end if;
	if (cc=68 and ll=321) then grbp<="011";
	end if;
	if (ll=321 and cc>=68 and cc<71) then grbp<="011";
	end if;
	if (ll=321 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=321 and cc>=136 and cc<138) then grbp<="011";
	end if;
	if (cc=147 and ll=321) then grbp<="011";
	end if;
	if (cc=209 and ll=321) then grbp<="011";
	end if;
	if (cc=33 and ll=322) then grbp<="011";
	end if;
	if (cc=56 and ll=322) then grbp<="011";
	end if;
	if (ll=322 and cc>=56 and cc<58) then grbp<="011";
	end if;
	if (cc=64 and ll=322) then grbp<="011";
	end if;
	if (cc=68 and ll=322) then grbp<="011";
	end if;
	if (cc=70 and ll=322) then grbp<="011";
	end if;
	if (cc=73 and ll=322) then grbp<="011";
	end if;
	if (cc=76 and ll=322) then grbp<="011";
	end if;
	if (cc=78 and ll=322) then grbp<="011";
	end if;
	if (cc=132 and ll=322) then grbp<="011";
	end if;
	if (cc=151 and ll=322) then grbp<="011";
	end if;
	if (cc=56 and ll=323) then grbp<="011";
	end if;
	if (ll=323 and cc>=56 and cc<58) then grbp<="011";
	end if;
	if (cc=65 and ll=323) then grbp<="011";
	end if;
	if (cc=67 and ll=323) then grbp<="011";
	end if;
	if (cc=69 and ll=323) then grbp<="011";
	end if;
	if (cc=73 and ll=323) then grbp<="011";
	end if;
	if (cc=79 and ll=323) then grbp<="011";
	end if;
	if (cc=32 and ll=324) then grbp<="011";
	end if;
	if (cc=56 and ll=324) then grbp<="011";
	end if;
	if (ll=324 and cc>=56 and cc<60) then grbp<="011";
	end if;
	if (cc=67 and ll=324) then grbp<="011";
	end if;
	if (cc=69 and ll=324) then grbp<="011";
	end if;
	if (cc=71 and ll=324) then grbp<="011";
	end if;
	if (cc=74 and ll=324) then grbp<="011";
	end if;
	if (cc=77 and ll=324) then grbp<="011";
	end if;
	if (cc=31 and ll=325) then grbp<="011";
	end if;
	if (cc=56 and ll=325) then grbp<="011";
	end if;
	if (ll=325 and cc>=56 and cc<59) then grbp<="011";
	end if;
	if (cc=65 and ll=325) then grbp<="011";
	end if;
	if (cc=71 and ll=325) then grbp<="011";
	end if;
	if (cc=73 and ll=325) then grbp<="011";
	end if;
	if (ll=325 and cc>=73 and cc<76) then grbp<="011";
	end if;
	if (cc=156 and ll=325) then grbp<="011";
	end if;
	if (cc=56 and ll=326) then grbp<="011";
	end if;
	if (ll=326 and cc>=56 and cc<61) then grbp<="011";
	end if;
	if (ll=326 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=71 and ll=326) then grbp<="011";
	end if;
	if (ll=326 and cc>=71 and cc<74) then grbp<="011";
	end if;
	if (cc=78 and ll=326) then grbp<="011";
	end if;
	if (cc=81 and ll=326) then grbp<="011";
	end if;
	if (cc=157 and ll=326) then grbp<="011";
	end if;
	if (cc=57 and ll=327) then grbp<="011";
	end if;
	if (ll=327 and cc>=57 and cc<59) then grbp<="011";
	end if;
	if (ll=327 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (ll=327 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=72 and ll=327) then grbp<="011";
	end if;
	if (ll=327 and cc>=72 and cc<74) then grbp<="011";
	end if;
	if (ll=327 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (ll=328 and cc>=57 and cc<59) then grbp<="011";
	end if;
	if (cc=65 and ll=328) then grbp<="011";
	end if;
	if (cc=73 and ll=328) then grbp<="011";
	end if;
	if (ll=328 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=328 and cc>=77 and cc<80) then grbp<="011";
	end if;
	if (cc=58 and ll=329) then grbp<="011";
	end if;
	if (ll=329 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (ll=329 and cc>=61 and cc<66) then grbp<="011";
	end if;
	if (cc=71 and ll=329) then grbp<="011";
	end if;
	if (cc=73 and ll=329) then grbp<="011";
	end if;
	if (ll=329 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (cc=79 and ll=329) then grbp<="011";
	end if;
	if (cc=81 and ll=329) then grbp<="011";
	end if;
	if (cc=59 and ll=330) then grbp<="011";
	end if;
	if (cc=63 and ll=330) then grbp<="011";
	end if;
	if (ll=330 and cc>=63 and cc<65) then grbp<="011";
	end if;
	if (cc=71 and ll=330) then grbp<="011";
	end if;
	if (ll=330 and cc>=71 and cc<78) then grbp<="011";
	end if;
	if (cc=162 and ll=330) then grbp<="011";
	end if;
	if (cc=34 and ll=331) then grbp<="011";
	end if;
	if (ll=331 and cc>=34 and cc<36) then grbp<="011";
	end if;
	if (ll=331 and cc>=58 and cc<61) then grbp<="011";
	end if;
	if (cc=70 and ll=331) then grbp<="011";
	end if;
	if (cc=72 and ll=331) then grbp<="011";
	end if;
	if (ll=331 and cc>=72 and cc<78) then grbp<="011";
	end if;
	if (cc=163 and ll=331) then grbp<="011";
	end if;
	if (cc=51 and ll=332) then grbp<="011";
	end if;
	if (cc=59 and ll=332) then grbp<="011";
	end if;
	if (ll=332 and cc>=59 and cc<62) then grbp<="011";
	end if;
	if (ll=332 and cc>=65 and cc<67) then grbp<="011";
	end if;
	if (cc=71 and ll=332) then grbp<="011";
	end if;
	if (ll=332 and cc>=71 and cc<77) then grbp<="011";
	end if;
	if (cc=0 and ll=333) then grbp<="011";
	end if;
	if (ll=333 and cc>=0 and cc<2) then grbp<="011";
	end if;
	if (cc=60 and ll=333) then grbp<="011";
	end if;
	if (ll=333 and cc>=60 and cc<64) then grbp<="011";
	end if;
	if (cc=68 and ll=333) then grbp<="011";
	end if;
	if (ll=333 and cc>=68 and cc<72) then grbp<="011";
	end if;
	if (ll=333 and cc>=73 and cc<78) then grbp<="011";
	end if;
	if (cc=82 and ll=333) then grbp<="011";
	end if;
	if (cc=84 and ll=333) then grbp<="011";
	end if;
	if (cc=165 and ll=333) then grbp<="011";
	end if;
	if (cc=0 and ll=334) then grbp<="011";
	end if;
	if (ll=334 and cc>=0 and cc<3) then grbp<="011";
	end if;
	if (cc=51 and ll=334) then grbp<="011";
	end if;
	if (cc=54 and ll=334) then grbp<="011";
	end if;
	if (cc=60 and ll=334) then grbp<="011";
	end if;
	if (ll=334 and cc>=60 and cc<65) then grbp<="011";
	end if;
	if (ll=334 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (ll=334 and cc>=73 and cc<78) then grbp<="011";
	end if;
	if (ll=335 and cc>=0 and cc<4) then grbp<="011";
	end if;
	if (cc=62 and ll=335) then grbp<="011";
	end if;
	if (ll=335 and cc>=62 and cc<64) then grbp<="011";
	end if;
	if (ll=335 and cc>=69 and cc<73) then grbp<="011";
	end if;
	if (ll=335 and cc>=75 and cc<78) then grbp<="011";
	end if;
	if (ll=336 and cc>=0 and cc<5) then grbp<="011";
	end if;
	if (ll=336 and cc>=44 and cc<47) then grbp<="011";
	end if;
	if (ll=336 and cc>=50 and cc<52) then grbp<="011";
	end if;
	if (ll=336 and cc>=62 and cc<65) then grbp<="011";
	end if;
	if (ll=336 and cc>=70 and cc<74) then grbp<="011";
	end if;
	if (ll=336 and cc>=75 and cc<78) then grbp<="011";
	end if;
	if (ll=337 and cc>=0 and cc<4) then grbp<="011";
	end if;
	if (cc=31 and ll=337) then grbp<="011";
	end if;
	if (cc=45 and ll=337) then grbp<="011";
	end if;
	if (ll=337 and cc>=45 and cc<51) then grbp<="011";
	end if;
	if (cc=62 and ll=337) then grbp<="011";
	end if;
	if (ll=337 and cc>=62 and cc<64) then grbp<="011";
	end if;
	if (ll=337 and cc>=70 and cc<74) then grbp<="011";
	end if;
	if (ll=337 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=168 and ll=337) then grbp<="011";
	end if;
	if (cc=0 and ll=338) then grbp<="011";
	end if;
	if (ll=338 and cc>=0 and cc<3) then grbp<="011";
	end if;
	if (ll=338 and cc>=5 and cc<7) then grbp<="011";
	end if;
	if (ll=338 and cc>=46 and cc<50) then grbp<="011";
	end if;
	if (ll=338 and cc>=57 and cc<59) then grbp<="011";
	end if;
	if (ll=338 and cc>=71 and cc<74) then grbp<="011";
	end if;
	if (ll=338 and cc>=75 and cc<79) then grbp<="011";
	end if;
	if (ll=339 and cc>=0 and cc<3) then grbp<="011";
	end if;
	if (cc=57 and ll=339) then grbp<="011";
	end if;
	if (cc=62 and ll=339) then grbp<="011";
	end if;
	if (cc=71 and ll=339) then grbp<="011";
	end if;
	if (ll=339 and cc>=71 and cc<76) then grbp<="011";
	end if;
	if (cc=82 and ll=339) then grbp<="011";
	end if;
	if (cc=1 and ll=340) then grbp<="011";
	end if;
	if (cc=7 and ll=340) then grbp<="011";
	end if;
	if (cc=55 and ll=340) then grbp<="011";
	end if;
	if (ll=340 and cc>=55 and cc<57) then grbp<="011";
	end if;
	if (ll=340 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=72 and ll=340) then grbp<="011";
	end if;
	if (ll=340 and cc>=72 and cc<76) then grbp<="011";
	end if;
	if (cc=1 and ll=341) then grbp<="011";
	end if;
	if (ll=341 and cc>=1 and cc<3) then grbp<="011";
	end if;
	if (ll=341 and cc>=7 and cc<9) then grbp<="011";
	end if;
	if (cc=61 and ll=341) then grbp<="011";
	end if;
	if (ll=341 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=341 and cc>=69 and cc<71) then grbp<="011";
	end if;
	if (ll=341 and cc>=72 and cc<76) then grbp<="011";
	end if;
	if (cc=83 and ll=341) then grbp<="011";
	end if;
	if (ll=341 and cc>=83 and cc<85) then grbp<="011";
	end if;
	if (cc=2 and ll=342) then grbp<="011";
	end if;
	if (cc=7 and ll=342) then grbp<="011";
	end if;
	if (ll=342 and cc>=7 and cc<9) then grbp<="011";
	end if;
	if (ll=342 and cc>=32 and cc<34) then grbp<="011";
	end if;
	if (ll=342 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=73 and ll=342) then grbp<="011";
	end if;
	if (cc=75 and ll=342) then grbp<="011";
	end if;
	if (ll=342 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (ll=342 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=2 and ll=343) then grbp<="011";
	end if;
	if (cc=9 and ll=343) then grbp<="011";
	end if;
	if (cc=62 and ll=343) then grbp<="011";
	end if;
	if (cc=70 and ll=343) then grbp<="011";
	end if;
	if (ll=343 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=343 and cc>=73 and cc<81) then grbp<="011";
	end if;
	if (cc=9 and ll=344) then grbp<="011";
	end if;
	if (cc=70 and ll=344) then grbp<="011";
	end if;
	if (ll=344 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=344 and cc>=73 and cc<81) then grbp<="011";
	end if;
	if (cc=3 and ll=345) then grbp<="011";
	end if;
	if (cc=9 and ll=345) then grbp<="011";
	end if;
	if (cc=63 and ll=345) then grbp<="011";
	end if;
	if (cc=71 and ll=345) then grbp<="011";
	end if;
	if (cc=75 and ll=345) then grbp<="011";
	end if;
	if (ll=345 and cc>=75 and cc<81) then grbp<="011";
	end if;
	if (ll=346 and cc>=3 and cc<5) then grbp<="011";
	end if;
	if (cc=71 and ll=346) then grbp<="011";
	end if;
	if (ll=346 and cc>=71 and cc<79) then grbp<="011";
	end if;
	if (cc=199 and ll=346) then grbp<="011";
	end if;
	if (cc=4 and ll=347) then grbp<="011";
	end if;
	if (cc=72 and ll=347) then grbp<="011";
	end if;
	if (ll=347 and cc>=72 and cc<79) then grbp<="011";
	end if;
	if (cc=85 and ll=347) then grbp<="011";
	end if;
	if (cc=173 and ll=347) then grbp<="011";
	end if;
	if (cc=4 and ll=348) then grbp<="011";
	end if;
	if (cc=51 and ll=348) then grbp<="011";
	end if;
	if (cc=59 and ll=348) then grbp<="011";
	end if;
	if (cc=65 and ll=348) then grbp<="011";
	end if;
	if (cc=73 and ll=348) then grbp<="011";
	end if;
	if (ll=348 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=348 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=85 and ll=348) then grbp<="011";
	end if;
	if (cc=4 and ll=349) then grbp<="011";
	end if;
	if (cc=51 and ll=349) then grbp<="011";
	end if;
	if (cc=68 and ll=349) then grbp<="011";
	end if;
	if (cc=73 and ll=349) then grbp<="011";
	end if;
	if (ll=349 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=349 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=85 and ll=349) then grbp<="011";
	end if;
	if (cc=4 and ll=350) then grbp<="011";
	end if;
	if (cc=32 and ll=350) then grbp<="011";
	end if;
	if (cc=51 and ll=350) then grbp<="011";
	end if;
	if (cc=66 and ll=350) then grbp<="011";
	end if;
	if (cc=68 and ll=350) then grbp<="011";
	end if;
	if (ll=350 and cc>=68 and cc<70) then grbp<="011";
	end if;
	if (ll=350 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=350 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=85 and ll=350) then grbp<="011";
	end if;
	if (cc=174 and ll=350) then grbp<="011";
	end if;
	if (cc=4 and ll=351) then grbp<="011";
	end if;
	if (cc=51 and ll=351) then grbp<="011";
	end if;
	if (cc=66 and ll=351) then grbp<="011";
	end if;
	if (cc=69 and ll=351) then grbp<="011";
	end if;
	if (ll=351 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (ll=351 and cc>=74 and cc<79) then grbp<="011";
	end if;
	if (cc=4 and ll=352) then grbp<="011";
	end if;
	if (cc=51 and ll=352) then grbp<="011";
	end if;
	if (cc=63 and ll=352) then grbp<="011";
	end if;
	if (cc=69 and ll=352) then grbp<="011";
	end if;
	if (ll=352 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=79 and ll=352) then grbp<="011";
	end if;
	if (cc=85 and ll=352) then grbp<="011";
	end if;
	if (ll=352 and cc>=85 and cc<87) then grbp<="011";
	end if;
	if (cc=51 and ll=353) then grbp<="011";
	end if;
	if (cc=63 and ll=353) then grbp<="011";
	end if;
	if (cc=69 and ll=353) then grbp<="011";
	end if;
	if (ll=353 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=80 and ll=353) then grbp<="011";
	end if;
	if (cc=33 and ll=354) then grbp<="011";
	end if;
	if (cc=51 and ll=354) then grbp<="011";
	end if;
	if (cc=69 and ll=354) then grbp<="011";
	end if;
	if (ll=354 and cc>=69 and cc<71) then grbp<="011";
	end if;
	if (cc=68 and ll=355) then grbp<="011";
	end if;
	if (cc=70 and ll=355) then grbp<="011";
	end if;
	if (cc=76 and ll=355) then grbp<="011";
	end if;
	if (cc=79 and ll=355) then grbp<="011";
	end if;
	if (cc=81 and ll=355) then grbp<="011";
	end if;
	if (cc=32 and ll=356) then grbp<="011";
	end if;
	if (cc=50 and ll=356) then grbp<="011";
	end if;
	if (ll=356 and cc>=50 and cc<52) then grbp<="011";
	end if;
	if (cc=68 and ll=356) then grbp<="011";
	end if;
	if (cc=70 and ll=356) then grbp<="011";
	end if;
	if (cc=76 and ll=356) then grbp<="011";
	end if;
	if (cc=78 and ll=356) then grbp<="011";
	end if;
	if (ll=356 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=50 and ll=357) then grbp<="011";
	end if;
	if (ll=357 and cc>=50 and cc<52) then grbp<="011";
	end if;
	if (ll=357 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (ll=357 and cc>=76 and cc<80) then grbp<="011";
	end if;
	if (ll=358 and cc>=50 and cc<52) then grbp<="011";
	end if;
	if (ll=358 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=358 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=50 and ll=359) then grbp<="011";
	end if;
	if (ll=359 and cc>=50 and cc<52) then grbp<="011";
	end if;
	if (ll=359 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=359 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=85 and ll=359) then grbp<="011";
	end if;
	if (cc=32 and ll=360) then grbp<="011";
	end if;
	if (cc=49 and ll=360) then grbp<="011";
	end if;
	if (ll=360 and cc>=49 and cc<52) then grbp<="011";
	end if;
	if (ll=360 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=360 and cc>=77 and cc<79) then grbp<="011";
	end if;
	if (cc=83 and ll=360) then grbp<="011";
	end if;
	if (ll=360 and cc>=83 and cc<85) then grbp<="011";
	end if;
	if (cc=49 and ll=361) then grbp<="011";
	end if;
	if (cc=70 and ll=361) then grbp<="011";
	end if;
	if (ll=361 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (ll=361 and cc>=77 and cc<79) then grbp<="011";
	end if;
	if (cc=82 and ll=361) then grbp<="011";
	end if;
	if (cc=84 and ll=361) then grbp<="011";
	end if;
	if (cc=87 and ll=361) then grbp<="011";
	end if;
	if (cc=5 and ll=362) then grbp<="011";
	end if;
	if (cc=48 and ll=362) then grbp<="011";
	end if;
	if (ll=362 and cc>=48 and cc<50) then grbp<="011";
	end if;
	if (ll=362 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (ll=362 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=84 and ll=362) then grbp<="011";
	end if;
	if (cc=87 and ll=362) then grbp<="011";
	end if;
	if (cc=5 and ll=363) then grbp<="011";
	end if;
	if (cc=48 and ll=363) then grbp<="011";
	end if;
	if (cc=71 and ll=363) then grbp<="011";
	end if;
	if (ll=363 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (ll=363 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (ll=363 and cc>=81 and cc<84) then grbp<="011";
	end if;
	if (cc=47 and ll=364) then grbp<="011";
	end if;
	if (cc=71 and ll=364) then grbp<="011";
	end if;
	if (ll=364 and cc>=71 and cc<78) then grbp<="011";
	end if;
	if (ll=364 and cc>=80 and cc<82) then grbp<="011";
	end if;
	if (cc=50 and ll=365) then grbp<="011";
	end if;
	if (cc=72 and ll=365) then grbp<="011";
	end if;
	if (ll=365 and cc>=72 and cc<78) then grbp<="011";
	end if;
	if (ll=365 and cc>=81 and cc<83) then grbp<="011";
	end if;
	if (cc=32 and ll=366) then grbp<="011";
	end if;
	if (cc=50 and ll=366) then grbp<="011";
	end if;
	if (cc=73 and ll=366) then grbp<="011";
	end if;
	if (ll=366 and cc>=73 and cc<80) then grbp<="011";
	end if;
	if (ll=366 and cc>=81 and cc<83) then grbp<="011";
	end if;
	if (cc=32 and ll=367) then grbp<="011";
	end if;
	if (cc=73 and ll=367) then grbp<="011";
	end if;
	if (ll=367 and cc>=73 and cc<80) then grbp<="011";
	end if;
	if (cc=87 and ll=367) then grbp<="011";
	end if;
	if (ll=367 and cc>=87 and cc<89) then grbp<="011";
	end if;
	if (cc=32 and ll=368) then grbp<="011";
	end if;
	if (cc=74 and ll=368) then grbp<="011";
	end if;
	if (cc=76 and ll=368) then grbp<="011";
	end if;
	if (ll=368 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (cc=88 and ll=368) then grbp<="011";
	end if;
	if (ll=368 and cc>=88 and cc<92) then grbp<="011";
	end if;
	if (cc=31 and ll=369) then grbp<="011";
	end if;
	if (ll=369 and cc>=31 and cc<33) then grbp<="011";
	end if;
	if (ll=369 and cc>=74 and cc<80) then grbp<="011";
	end if;
	if (ll=369 and cc>=90 and cc<96) then grbp<="011";
	end if;
	if (cc=74 and ll=370) then grbp<="011";
	end if;
	if (ll=370 and cc>=74 and cc<80) then grbp<="011";
	end if;
	if (cc=11 and ll=371) then grbp<="011";
	end if;
	if (cc=31 and ll=371) then grbp<="011";
	end if;
	if (cc=67 and ll=371) then grbp<="011";
	end if;
	if (cc=74 and ll=371) then grbp<="011";
	end if;
	if (cc=76 and ll=371) then grbp<="011";
	end if;
	if (ll=371 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=81 and ll=371) then grbp<="011";
	end if;
	if (cc=84 and ll=371) then grbp<="011";
	end if;
	if (cc=96 and ll=371) then grbp<="011";
	end if;
	if (cc=11 and ll=372) then grbp<="011";
	end if;
	if (cc=74 and ll=372) then grbp<="011";
	end if;
	if (ll=372 and cc>=74 and cc<82) then grbp<="011";
	end if;
	if (ll=373 and cc>=74 and cc<82) then grbp<="011";
	end if;
	if (ll=374 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=82 and ll=374) then grbp<="011";
	end if;
	if (cc=188 and ll=374) then grbp<="011";
	end if;
	if (cc=11 and ll=375) then grbp<="011";
	end if;
	if (cc=66 and ll=375) then grbp<="011";
	end if;
	if (cc=69 and ll=375) then grbp<="011";
	end if;
	if (cc=72 and ll=375) then grbp<="011";
	end if;
	if (cc=77 and ll=375) then grbp<="011";
	end if;
	if (cc=81 and ll=375) then grbp<="011";
	end if;
	if (cc=72 and ll=376) then grbp<="011";
	end if;
	if (ll=376 and cc>=72 and cc<78) then grbp<="011";
	end if;
	if (ll=376 and cc>=81 and cc<84) then grbp<="011";
	end if;
	if (ll=377 and cc>=75 and cc<79) then grbp<="011";
	end if;
	if (ll=377 and cc>=82 and cc<85) then grbp<="011";
	end if;
	if (cc=6 and ll=378) then grbp<="011";
	end if;
	if (cc=73 and ll=378) then grbp<="011";
	end if;
	if (ll=378 and cc>=73 and cc<78) then grbp<="011";
	end if;
	if (cc=84 and ll=378) then grbp<="011";
	end if;
	if (cc=6 and ll=379) then grbp<="011";
	end if;
	if (cc=76 and ll=379) then grbp<="011";
	end if;
	if (ll=379 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (ll=379 and cc>=82 and cc<84) then grbp<="011";
	end if;
	if (cc=6 and ll=380) then grbp<="011";
	end if;
	if (cc=70 and ll=380) then grbp<="011";
	end if;
	if (cc=78 and ll=380) then grbp<="011";
	end if;
	if (cc=83 and ll=380) then grbp<="011";
	end if;
	if (cc=32 and ll=381) then grbp<="011";
	end if;
	if (cc=70 and ll=381) then grbp<="011";
	end if;
	if (cc=83 and ll=381) then grbp<="011";
	end if;
	if (cc=6 and ll=382) then grbp<="011";
	end if;
	if (cc=32 and ll=382) then grbp<="011";
	end if;
	if (cc=69 and ll=382) then grbp<="011";
	end if;
	if (ll=382 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=6 and ll=383) then grbp<="011";
	end if;
	if (cc=69 and ll=383) then grbp<="011";
	end if;
	if (ll=383 and cc>=69 and cc<72) then grbp<="011";
	end if;
	if (cc=85 and ll=383) then grbp<="011";
	end if;
	if (cc=6 and ll=384) then grbp<="011";
	end if;
	if (cc=70 and ll=384) then grbp<="011";
	end if;
	if (ll=384 and cc>=70 and cc<72) then grbp<="011";
	end if;
	if (cc=85 and ll=384) then grbp<="011";
	end if;
	if (cc=67 and ll=385) then grbp<="011";
	end if;
	if (cc=70 and ll=385) then grbp<="011";
	end if;
	if (ll=385 and cc>=70 and cc<73) then grbp<="011";
	end if;
	if (cc=68 and ll=386) then grbp<="011";
	end if;
	if (ll=386 and cc>=68 and cc<72) then grbp<="011";
	end if;
	if (cc=68 and ll=387) then grbp<="011";
	end if;
	if (ll=387 and cc>=68 and cc<72) then grbp<="011";
	end if;
	if (cc=81 and ll=387) then grbp<="011";
	end if;
	if (cc=6 and ll=388) then grbp<="011";
	end if;
	if (cc=71 and ll=388) then grbp<="011";
	end if;
	if (ll=388 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (cc=6 and ll=389) then grbp<="011";
	end if;
	if (cc=71 and ll=389) then grbp<="011";
	end if;
	if (ll=389 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (cc=77 and ll=389) then grbp<="011";
	end if;
	if (cc=79 and ll=389) then grbp<="011";
	end if;
	if (cc=71 and ll=390) then grbp<="011";
	end if;
	if (ll=390 and cc>=71 and cc<74) then grbp<="011";
	end if;
	if (cc=79 and ll=390) then grbp<="011";
	end if;
	if (cc=70 and ll=391) then grbp<="011";
	end if;
	if (ll=391 and cc>=70 and cc<76) then grbp<="011";
	end if;
	if (ll=392 and cc>=71 and cc<73) then grbp<="011";
	end if;
	if (ll=392 and cc>=74 and cc<78) then grbp<="011";
	end if;
	if (cc=75 and ll=393) then grbp<="011";
	end if;
	if (ll=393 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (ll=393 and cc>=79 and cc<81) then grbp<="011";
	end if;
	if (cc=75 and ll=394) then grbp<="011";
	end if;
	if (ll=394 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (ll=394 and cc>=79 and cc<81) then grbp<="011";
	end if;
	if (ll=395 and cc>=73 and cc<75) then grbp<="011";
	end if;
	if (ll=395 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=74 and ll=396) then grbp<="011";
	end if;
	if (ll=396 and cc>=74 and cc<76) then grbp<="011";
	end if;
	if (ll=396 and cc>=77 and cc<80) then grbp<="011";
	end if;
	if (cc=74 and ll=397) then grbp<="011";
	end if;
	if (ll=397 and cc>=74 and cc<76) then grbp<="011";
	end if;
	if (cc=80 and ll=397) then grbp<="011";
	end if;
	if (ll=397 and cc>=80 and cc<82) then grbp<="011";
	end if;
	if (ll=398 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (ll=399 and cc>=78 and cc<80) then grbp<="011";
	end if;
	if (cc=78 and ll=400) then grbp<="011";
	end if;
	if (ll=400 and cc>=78 and cc<81) then grbp<="011";
	end if;
	if (cc=75 and ll=401) then grbp<="011";
	end if;
	if (ll=401 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (ll=401 and cc>=79 and cc<81) then grbp<="011";
	end if;
	if (cc=75 and ll=402) then grbp<="011";
	end if;
	if (ll=402 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (cc=77 and ll=403) then grbp<="011";
	end if;
	if (cc=76 and ll=404) then grbp<="011";
	end if;
	if (ll=404 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=227 and ll=404) then grbp<="011";
	end if;
	if (cc=7 and ll=405) then grbp<="011";
	end if;
	if (cc=54 and ll=405) then grbp<="011";
	end if;
	if (cc=70 and ll=405) then grbp<="011";
	end if;
	if (cc=76 and ll=405) then grbp<="011";
	end if;
	if (ll=405 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=212 and ll=405) then grbp<="011";
	end if;
	if (cc=218 and ll=405) then grbp<="011";
	end if;
	if (cc=244 and ll=405) then grbp<="011";
	end if;
	if (cc=7 and ll=406) then grbp<="011";
	end if;
	if (cc=54 and ll=406) then grbp<="011";
	end if;
	if (cc=70 and ll=406) then grbp<="011";
	end if;
	if (cc=76 and ll=406) then grbp<="011";
	end if;
	if (cc=78 and ll=406) then grbp<="011";
	end if;
	if (cc=205 and ll=406) then grbp<="011";
	end if;
	if (cc=218 and ll=406) then grbp<="011";
	end if;
	if (cc=223 and ll=406) then grbp<="011";
	end if;
	if (ll=406 and cc>=223 and cc<226) then grbp<="011";
	end if;
	if (cc=59 and ll=407) then grbp<="011";
	end if;
	if (cc=70 and ll=407) then grbp<="011";
	end if;
	if (cc=75 and ll=407) then grbp<="011";
	end if;
	if (ll=407 and cc>=75 and cc<77) then grbp<="011";
	end if;
	if (cc=191 and ll=407) then grbp<="011";
	end if;
	if (cc=216 and ll=407) then grbp<="011";
	end if;
	if (cc=218 and ll=407) then grbp<="011";
	end if;
	if (cc=225 and ll=407) then grbp<="011";
	end if;
	if (cc=230 and ll=407) then grbp<="011";
	end if;
	if (cc=235 and ll=407) then grbp<="011";
	end if;
	if (cc=7 and ll=408) then grbp<="011";
	end if;
	if (cc=59 and ll=408) then grbp<="011";
	end if;
	if (cc=71 and ll=408) then grbp<="011";
	end if;
	if (cc=75 and ll=408) then grbp<="011";
	end if;
	if (ll=408 and cc>=75 and cc<78) then grbp<="011";
	end if;
	if (cc=218 and ll=408) then grbp<="011";
	end if;
	if (cc=230 and ll=408) then grbp<="011";
	end if;
	if (cc=7 and ll=409) then grbp<="011";
	end if;
	if (cc=59 and ll=409) then grbp<="011";
	end if;
	if (cc=71 and ll=409) then grbp<="011";
	end if;
	if (cc=75 and ll=409) then grbp<="011";
	end if;
	if (ll=409 and cc>=75 and cc<80) then grbp<="011";
	end if;
	if (cc=200 and ll=409) then grbp<="011";
	end if;
	if (cc=218 and ll=409) then grbp<="011";
	end if;
	if (cc=230 and ll=409) then grbp<="011";
	end if;
	if (cc=59 and ll=410) then grbp<="011";
	end if;
	if (ll=410 and cc>=59 and cc<62) then grbp<="011";
	end if;
	if (ll=410 and cc>=75 and cc<78) then grbp<="011";
	end if;
	if (cc=190 and ll=410) then grbp<="011";
	end if;
	if (cc=196 and ll=410) then grbp<="011";
	end if;
	if (cc=230 and ll=410) then grbp<="011";
	end if;
	if (cc=237 and ll=410) then grbp<="011";
	end if;
	if (cc=240 and ll=410) then grbp<="011";
	end if;
	if (ll=410 and cc>=240 and cc<242) then grbp<="011";
	end if;
	if (ll=411 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (cc=76 and ll=411) then grbp<="011";
	end if;
	if (ll=411 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (ll=411 and cc>=79 and cc<81) then grbp<="011";
	end if;
	if (cc=230 and ll=411) then grbp<="011";
	end if;
	if (cc=237 and ll=411) then grbp<="011";
	end if;
	if (ll=411 and cc>=237 and cc<239) then grbp<="011";
	end if;
	if (cc=60 and ll=412) then grbp<="011";
	end if;
	if (ll=412 and cc>=60 and cc<62) then grbp<="011";
	end if;
	if (cc=76 and ll=412) then grbp<="011";
	end if;
	if (ll=412 and cc>=76 and cc<78) then grbp<="011";
	end if;
	if (cc=220 and ll=412) then grbp<="011";
	end if;
	if (cc=226 and ll=412) then grbp<="011";
	end if;
	if (cc=230 and ll=412) then grbp<="011";
	end if;
	if (cc=243 and ll=412) then grbp<="011";
	end if;
	if (cc=59 and ll=413) then grbp<="011";
	end if;
	if (cc=61 and ll=413) then grbp<="011";
	end if;
	if (cc=67 and ll=413) then grbp<="011";
	end if;
	if (cc=76 and ll=413) then grbp<="011";
	end if;
	if (ll=413 and cc>=76 and cc<79) then grbp<="011";
	end if;
	if (ll=413 and cc>=195 and cc<197) then grbp<="011";
	end if;
	if (cc=208 and ll=413) then grbp<="011";
	end if;
	if (cc=221 and ll=413) then grbp<="011";
	end if;
	if (cc=234 and ll=413) then grbp<="011";
	end if;
	if (cc=238 and ll=413) then grbp<="011";
	end if;
	if (cc=59 and ll=414) then grbp<="011";
	end if;
	if (cc=61 and ll=414) then grbp<="011";
	end if;
	if (ll=414 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=414 and cc>=66 and cc<68) then grbp<="011";
	end if;
	if (cc=77 and ll=414) then grbp<="011";
	end if;
	if (ll=414 and cc>=77 and cc<79) then grbp<="011";
	end if;
	if (cc=59 and ll=415) then grbp<="011";
	end if;
	if (cc=61 and ll=415) then grbp<="011";
	end if;
	if (ll=415 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (ll=415 and cc>=66 and cc<68) then grbp<="011";
	end if;
	if (cc=78 and ll=415) then grbp<="011";
	end if;
	if (cc=53 and ll=416) then grbp<="011";
	end if;
	if (cc=58 and ll=416) then grbp<="011";
	end if;
	if (ll=416 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (ll=416 and cc>=61 and cc<63) then grbp<="011";
	end if;
	if (cc=79 and ll=416) then grbp<="011";
	end if;
	if (cc=186 and ll=416) then grbp<="011";
	end if;
	if (cc=53 and ll=417) then grbp<="011";
	end if;
	if (cc=58 and ll=417) then grbp<="011";
	end if;
	if (ll=417 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (cc=74 and ll=417) then grbp<="011";
	end if;
	if (cc=53 and ll=418) then grbp<="011";
	end if;
	if (cc=58 and ll=418) then grbp<="011";
	end if;
	if (ll=418 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (ll=418 and cc>=62 and cc<64) then grbp<="011";
	end if;
	if (cc=79 and ll=418) then grbp<="011";
	end if;
	if (cc=81 and ll=418) then grbp<="011";
	end if;
	if (cc=53 and ll=419) then grbp<="011";
	end if;
	if (cc=58 and ll=419) then grbp<="011";
	end if;
	if (ll=419 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (cc=68 and ll=419) then grbp<="011";
	end if;
	if (cc=79 and ll=419) then grbp<="011";
	end if;
	if (cc=81 and ll=419) then grbp<="011";
	end if;
	if (cc=59 and ll=420) then grbp<="011";
	end if;
	if (cc=79 and ll=420) then grbp<="011";
	end if;
	if (cc=81 and ll=420) then grbp<="011";
	end if;
	if (ll=420 and cc>=81 and cc<83) then grbp<="011";
	end if;
	if (cc=59 and ll=421) then grbp<="011";
	end if;
	if (cc=63 and ll=421) then grbp<="011";
	end if;
	if (ll=421 and cc>=63 and cc<65) then grbp<="011";
	end if;
	if (ll=421 and cc>=82 and cc<84) then grbp<="011";
	end if;
	if (cc=58 and ll=422) then grbp<="011";
	end if;
	if (ll=422 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (cc=68 and ll=422) then grbp<="011";
	end if;
	if (cc=82 and ll=422) then grbp<="011";
	end if;
	if (cc=58 and ll=423) then grbp<="011";
	end if;
	if (ll=423 and cc>=58 and cc<60) then grbp<="011";
	end if;
	if (ll=423 and cc>=64 and cc<66) then grbp<="011";
	end if;
	if (cc=84 and ll=423) then grbp<="011";
	end if;
	if (cc=59 and ll=424) then grbp<="011";
	end if;
	if (cc=64 and ll=424) then grbp<="011";
	end if;
	if (ll=424 and cc>=64 and cc<66) then grbp<="011";
	end if;
	if (cc=80 and ll=424) then grbp<="011";
	end if;
	if (cc=84 and ll=424) then grbp<="011";
	end if;
	if (cc=188 and ll=424) then grbp<="011";
	end if;


	if (cc=1 and ll=0) then grbp<="111";
	end if;
	if (cc=198 and ll=0) then grbp<="111";
	end if;
	if (ll=0 and cc>=198 and cc<206) then grbp<="111";
	end if;
	if (cc=1 and ll=1) then grbp<="111";
	end if;
	if (cc=198 and ll=1) then grbp<="111";
	end if;
	if (ll=1 and cc>=198 and cc<206) then grbp<="111";
	end if;
	if (cc=1 and ll=2) then grbp<="111";
	end if;
	if (cc=198 and ll=2) then grbp<="111";
	end if;
	if (ll=2 and cc>=198 and cc<206) then grbp<="111";
	end if;
	if (cc=1 and ll=3) then grbp<="111";
	end if;
	if (cc=198 and ll=3) then grbp<="111";
	end if;
	if (ll=3 and cc>=198 and cc<206) then grbp<="111";
	end if;
	if (cc=199 and ll=4) then grbp<="111";
	end if;
	if (ll=4 and cc>=199 and cc<207) then grbp<="111";
	end if;
	if (ll=5 and cc>=199 and cc<207) then grbp<="111";
	end if;
	if (ll=6 and cc>=199 and cc<207) then grbp<="111";
	end if;
	if (ll=7 and cc>=200 and cc<207) then grbp<="111";
	end if;
	if (ll=8 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=9 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=10 and cc>=201 and cc<209) then grbp<="111";
	end if;
	if (ll=11 and cc>=201 and cc<209) then grbp<="111";
	end if;
	if (ll=12 and cc>=202 and cc<210) then grbp<="111";
	end if;
	if (ll=13 and cc>=201 and cc<210) then grbp<="111";
	end if;
	if (ll=14 and cc>=202 and cc<210) then grbp<="111";
	end if;
	if (ll=15 and cc>=202 and cc<210) then grbp<="111";
	end if;
	if (ll=16 and cc>=203 and cc<211) then grbp<="111";
	end if;
	if (ll=17 and cc>=203 and cc<211) then grbp<="111";
	end if;
	if (ll=18 and cc>=203 and cc<211) then grbp<="111";
	end if;
	if (ll=19 and cc>=204 and cc<212) then grbp<="111";
	end if;
	if (ll=20 and cc>=204 and cc<212) then grbp<="111";
	end if;
	if (ll=21 and cc>=204 and cc<213) then grbp<="111";
	end if;
	if (ll=22 and cc>=205 and cc<213) then grbp<="111";
	end if;
	if (ll=23 and cc>=205 and cc<213) then grbp<="111";
	end if;
	if (ll=24 and cc>=206 and cc<213) then grbp<="111";
	end if;
	if (ll=25 and cc>=206 and cc<214) then grbp<="111";
	end if;
	if (ll=26 and cc>=208 and cc<215) then grbp<="111";
	end if;
	if (ll=27 and cc>=208 and cc<215) then grbp<="111";
	end if;
	if (ll=28 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (ll=29 and cc>=207 and cc<216) then grbp<="111";
	end if;
	if (ll=30 and cc>=207 and cc<216) then grbp<="111";
	end if;
	if (ll=31 and cc>=208 and cc<216) then grbp<="111";
	end if;
	if (ll=32 and cc>=208 and cc<216) then grbp<="111";
	end if;
	if (ll=33 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=34 and cc>=209 and cc<217) then grbp<="111";
	end if;
	if (ll=35 and cc>=209 and cc<217) then grbp<="111";
	end if;
	if (ll=36 and cc>=209 and cc<218) then grbp<="111";
	end if;
	if (cc=111 and ll=37) then grbp<="111";
	end if;
	if (cc=113 and ll=37) then grbp<="111";
	end if;
	if (cc=210 and ll=37) then grbp<="111";
	end if;
	if (ll=37 and cc>=210 and cc<218) then grbp<="111";
	end if;
	if (ll=38 and cc>=108 and cc<118) then grbp<="111";
	end if;
	if (ll=38 and cc>=210 and cc<218) then grbp<="111";
	end if;
	if (cc=102 and ll=39) then grbp<="111";
	end if;
	if (cc=106 and ll=39) then grbp<="111";
	end if;
	if (ll=39 and cc>=106 and cc<119) then grbp<="111";
	end if;
	if (ll=39 and cc>=210 and cc<219) then grbp<="111";
	end if;
	if (ll=40 and cc>=105 and cc<121) then grbp<="111";
	end if;
	if (ll=40 and cc>=211 and cc<219) then grbp<="111";
	end if;
	if (ll=41 and cc>=99 and cc<102) then grbp<="111";
	end if;
	if (ll=41 and cc>=104 and cc<123) then grbp<="111";
	end if;
	if (ll=41 and cc>=211 and cc<220) then grbp<="111";
	end if;
	if (cc=99 and ll=42) then grbp<="111";
	end if;
	if (cc=101 and ll=42) then grbp<="111";
	end if;
	if (ll=42 and cc>=101 and cc<125) then grbp<="111";
	end if;
	if (ll=42 and cc>=211 and cc<220) then grbp<="111";
	end if;
	if (ll=43 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=43 and cc>=100 and cc<102) then grbp<="111";
	end if;
	if (ll=43 and cc>=103 and cc<126) then grbp<="111";
	end if;
	if (ll=43 and cc>=212 and cc<220) then grbp<="111";
	end if;
	if (cc=103 and ll=44) then grbp<="111";
	end if;
	if (ll=44 and cc>=103 and cc<128) then grbp<="111";
	end if;
	if (ll=44 and cc>=212 and cc<221) then grbp<="111";
	end if;
	if (cc=101 and ll=45) then grbp<="111";
	end if;
	if (ll=45 and cc>=101 and cc<103) then grbp<="111";
	end if;
	if (ll=45 and cc>=104 and cc<129) then grbp<="111";
	end if;
	if (ll=45 and cc>=213 and cc<221) then grbp<="111";
	end if;
	if (cc=101 and ll=46) then grbp<="111";
	end if;
	if (cc=103 and ll=46) then grbp<="111";
	end if;
	if (ll=46 and cc>=103 and cc<130) then grbp<="111";
	end if;
	if (ll=46 and cc>=213 and cc<222) then grbp<="111";
	end if;
	if (cc=100 and ll=47) then grbp<="111";
	end if;
	if (cc=104 and ll=47) then grbp<="111";
	end if;
	if (ll=47 and cc>=104 and cc<131) then grbp<="111";
	end if;
	if (ll=47 and cc>=213 and cc<222) then grbp<="111";
	end if;
	if (cc=101 and ll=48) then grbp<="111";
	end if;
	if (cc=103 and ll=48) then grbp<="111";
	end if;
	if (cc=105 and ll=48) then grbp<="111";
	end if;
	if (ll=48 and cc>=105 and cc<131) then grbp<="111";
	end if;
	if (ll=48 and cc>=213 and cc<222) then grbp<="111";
	end if;
	if (cc=99 and ll=49) then grbp<="111";
	end if;
	if (cc=101 and ll=49) then grbp<="111";
	end if;
	if (cc=104 and ll=49) then grbp<="111";
	end if;
	if (ll=49 and cc>=104 and cc<132) then grbp<="111";
	end if;
	if (ll=49 and cc>=214 and cc<222) then grbp<="111";
	end if;
	if (cc=101 and ll=50) then grbp<="111";
	end if;
	if (cc=103 and ll=50) then grbp<="111";
	end if;
	if (cc=105 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=105 and cc<133) then grbp<="111";
	end if;
	if (ll=50 and cc>=214 and cc<222) then grbp<="111";
	end if;
	if (ll=51 and cc>=103 and cc<105) then grbp<="111";
	end if;
	if (ll=51 and cc>=106 and cc<134) then grbp<="111";
	end if;
	if (ll=51 and cc>=214 and cc<222) then grbp<="111";
	end if;
	if (cc=103 and ll=52) then grbp<="111";
	end if;
	if (cc=105 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=105 and cc<109) then grbp<="111";
	end if;
	if (ll=52 and cc>=110 and cc<135) then grbp<="111";
	end if;
	if (ll=52 and cc>=215 and cc<221) then grbp<="111";
	end if;
	if (cc=105 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=105 and cc<109) then grbp<="111";
	end if;
	if (cc=112 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=112 and cc<136) then grbp<="111";
	end if;
	if (ll=53 and cc>=215 and cc<221) then grbp<="111";
	end if;
	if (cc=105 and ll=54) then grbp<="111";
	end if;
	if (cc=107 and ll=54) then grbp<="111";
	end if;
	if (cc=109 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=109 and cc<137) then grbp<="111";
	end if;
	if (ll=54 and cc>=216 and cc<220) then grbp<="111";
	end if;
	if (cc=105 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=105 and cc<107) then grbp<="111";
	end if;
	if (ll=55 and cc>=108 and cc<137) then grbp<="111";
	end if;
	if (ll=55 and cc>=216 and cc<220) then grbp<="111";
	end if;
	if (ll=56 and cc>=107 and cc<138) then grbp<="111";
	end if;
	if (ll=56 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=57 and cc>=107 and cc<109) then grbp<="111";
	end if;
	if (ll=57 and cc>=110 and cc<139) then grbp<="111";
	end if;
	if (ll=57 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=58 and cc>=107 and cc<140) then grbp<="111";
	end if;
	if (cc=106 and ll=59) then grbp<="111";
	end if;
	if (cc=108 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=108 and cc<141) then grbp<="111";
	end if;
	if (ll=60 and cc>=108 and cc<141) then grbp<="111";
	end if;
	if (cc=109 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=109 and cc<142) then grbp<="111";
	end if;
	if (cc=110 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=110 and cc<144) then grbp<="111";
	end if;
	if (cc=110 and ll=63) then grbp<="111";
	end if;
	if (cc=112 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=112 and cc<145) then grbp<="111";
	end if;
	if (ll=64 and cc>=109 and cc<146) then grbp<="111";
	end if;
	if (cc=110 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=110 and cc<146) then grbp<="111";
	end if;
	if (cc=109 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=109 and cc<111) then grbp<="111";
	end if;
	if (ll=66 and cc>=112 and cc<146) then grbp<="111";
	end if;
	if (cc=111 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=111 and cc<147) then grbp<="111";
	end if;
	if (ll=68 and cc>=110 and cc<147) then grbp<="111";
	end if;
	if (ll=69 and cc>=111 and cc<148) then grbp<="111";
	end if;
	if (ll=70 and cc>=109 and cc<148) then grbp<="111";
	end if;
	if (cc=111 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=111 and cc<148) then grbp<="111";
	end if;
	if (ll=72 and cc>=109 and cc<149) then grbp<="111";
	end if;
	if (ll=73 and cc>=111 and cc<149) then grbp<="111";
	end if;
	if (cc=110 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=110 and cc<150) then grbp<="111";
	end if;
	if (cc=113 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=113 and cc<150) then grbp<="111";
	end if;
	if (ll=76 and cc>=111 and cc<151) then grbp<="111";
	end if;
	if (ll=77 and cc>=111 and cc<118) then grbp<="111";
	end if;
	if (ll=77 and cc>=119 and cc<151) then grbp<="111";
	end if;
	if (ll=78 and cc>=111 and cc<118) then grbp<="111";
	end if;
	if (ll=78 and cc>=119 and cc<151) then grbp<="111";
	end if;
	if (ll=79 and cc>=111 and cc<115) then grbp<="111";
	end if;
	if (ll=79 and cc>=118 and cc<152) then grbp<="111";
	end if;
	if (cc=109 and ll=80) then grbp<="111";
	end if;
	if (cc=111 and ll=80) then grbp<="111";
	end if;
	if (ll=80 and cc>=111 and cc<114) then grbp<="111";
	end if;
	if (ll=80 and cc>=117 and cc<153) then grbp<="111";
	end if;
	if (ll=81 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (ll=81 and cc>=116 and cc<154) then grbp<="111";
	end if;
	if (ll=82 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (ll=82 and cc>=115 and cc<155) then grbp<="111";
	end if;
	if (ll=82 and cc>=248 and cc<251) then grbp<="111";
	end if;
	if (ll=83 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (ll=83 and cc>=114 and cc<155) then grbp<="111";
	end if;
	if (cc=249 and ll=83) then grbp<="111";
	end if;
	if (cc=111 and ll=84) then grbp<="111";
	end if;
	if (cc=114 and ll=84) then grbp<="111";
	end if;
	if (ll=84 and cc>=114 and cc<156) then grbp<="111";
	end if;
	if (cc=248 and ll=84) then grbp<="111";
	end if;
	if (cc=113 and ll=85) then grbp<="111";
	end if;
	if (ll=85 and cc>=113 and cc<156) then grbp<="111";
	end if;
	if (ll=85 and cc>=247 and cc<250) then grbp<="111";
	end if;
	if (ll=86 and cc>=112 and cc<157) then grbp<="111";
	end if;
	if (ll=86 and cc>=247 and cc<250) then grbp<="111";
	end if;
	if (ll=87 and cc>=111 and cc<157) then grbp<="111";
	end if;
	if (ll=87 and cc>=245 and cc<249) then grbp<="111";
	end if;
	if (cc=64 and ll=88) then grbp<="111";
	end if;
	if (cc=110 and ll=88) then grbp<="111";
	end if;
	if (ll=88 and cc>=110 and cc<158) then grbp<="111";
	end if;
	if (cc=245 and ll=88) then grbp<="111";
	end if;
	if (ll=88 and cc>=245 and cc<247) then grbp<="111";
	end if;
	if (cc=64 and ll=89) then grbp<="111";
	end if;
	if (cc=109 and ll=89) then grbp<="111";
	end if;
	if (ll=89 and cc>=109 and cc<158) then grbp<="111";
	end if;
	if (cc=64 and ll=90) then grbp<="111";
	end if;
	if (cc=109 and ll=90) then grbp<="111";
	end if;
	if (ll=90 and cc>=109 and cc<158) then grbp<="111";
	end if;
	if (cc=245 and ll=90) then grbp<="111";
	end if;
	if (cc=249 and ll=90) then grbp<="111";
	end if;
	if (cc=64 and ll=91) then grbp<="111";
	end if;
	if (cc=108 and ll=91) then grbp<="111";
	end if;
	if (ll=91 and cc>=108 and cc<159) then grbp<="111";
	end if;
	if (ll=92 and cc>=107 and cc<159) then grbp<="111";
	end if;
	if (ll=92 and cc>=194 and cc<199) then grbp<="111";
	end if;
	if (cc=236 and ll=92) then grbp<="111";
	end if;
	if (cc=242 and ll=92) then grbp<="111";
	end if;
	if (cc=244 and ll=92) then grbp<="111";
	end if;
	if (cc=246 and ll=92) then grbp<="111";
	end if;
	if (ll=92 and cc>=246 and cc<249) then grbp<="111";
	end if;
	if (cc=106 and ll=93) then grbp<="111";
	end if;
	if (ll=93 and cc>=106 and cc<160) then grbp<="111";
	end if;
	if (ll=93 and cc>=194 and cc<202) then grbp<="111";
	end if;
	if (cc=244 and ll=93) then grbp<="111";
	end if;
	if (ll=93 and cc>=244 and cc<246) then grbp<="111";
	end if;
	if (cc=106 and ll=94) then grbp<="111";
	end if;
	if (ll=94 and cc>=106 and cc<160) then grbp<="111";
	end if;
	if (ll=94 and cc>=193 and cc<203) then grbp<="111";
	end if;
	if (ll=94 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (cc=63 and ll=95) then grbp<="111";
	end if;
	if (cc=105 and ll=95) then grbp<="111";
	end if;
	if (cc=107 and ll=95) then grbp<="111";
	end if;
	if (ll=95 and cc>=107 and cc<160) then grbp<="111";
	end if;
	if (ll=95 and cc>=192 and cc<204) then grbp<="111";
	end if;
	if (ll=95 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (ll=96 and cc>=62 and cc<64) then grbp<="111";
	end if;
	if (ll=96 and cc>=104 and cc<160) then grbp<="111";
	end if;
	if (ll=96 and cc>=191 and cc<204) then grbp<="111";
	end if;
	if (ll=96 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (ll=97 and cc>=62 and cc<64) then grbp<="111";
	end if;
	if (ll=97 and cc>=103 and cc<160) then grbp<="111";
	end if;
	if (ll=97 and cc>=190 and cc<204) then grbp<="111";
	end if;
	if (ll=97 and cc>=241 and cc<245) then grbp<="111";
	end if;
	if (cc=102 and ll=98) then grbp<="111";
	end if;
	if (ll=98 and cc>=102 and cc<161) then grbp<="111";
	end if;
	if (ll=98 and cc>=190 and cc<204) then grbp<="111";
	end if;
	if (ll=98 and cc>=240 and cc<243) then grbp<="111";
	end if;
	if (cc=62 and ll=99) then grbp<="111";
	end if;
	if (cc=101 and ll=99) then grbp<="111";
	end if;
	if (ll=99 and cc>=101 and cc<161) then grbp<="111";
	end if;
	if (ll=99 and cc>=189 and cc<204) then grbp<="111";
	end if;
	if (cc=238 and ll=99) then grbp<="111";
	end if;
	if (cc=240 and ll=99) then grbp<="111";
	end if;
	if (ll=99 and cc>=240 and cc<243) then grbp<="111";
	end if;
	if (ll=99 and cc>=245 and cc<247) then grbp<="111";
	end if;
	if (cc=101 and ll=100) then grbp<="111";
	end if;
	if (ll=100 and cc>=101 and cc<161) then grbp<="111";
	end if;
	if (ll=100 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=240 and ll=100) then grbp<="111";
	end if;
	if (ll=100 and cc>=240 and cc<242) then grbp<="111";
	end if;
	if (cc=245 and ll=100) then grbp<="111";
	end if;
	if (ll=100 and cc>=245 and cc<247) then grbp<="111";
	end if;
	if (cc=100 and ll=101) then grbp<="111";
	end if;
	if (ll=101 and cc>=100 and cc<107) then grbp<="111";
	end if;
	if (ll=101 and cc>=108 and cc<162) then grbp<="111";
	end if;
	if (ll=101 and cc>=187 and cc<205) then grbp<="111";
	end if;
	if (cc=243 and ll=101) then grbp<="111";
	end if;
	if (cc=246 and ll=101) then grbp<="111";
	end if;
	if (cc=61 and ll=102) then grbp<="111";
	end if;
	if (ll=102 and cc>=61 and cc<63) then grbp<="111";
	end if;
	if (ll=102 and cc>=99 and cc<162) then grbp<="111";
	end if;
	if (ll=102 and cc>=187 and cc<205) then grbp<="111";
	end if;
	if (ll=102 and cc>=237 and cc<243) then grbp<="111";
	end if;
	if (ll=103 and cc>=61 and cc<63) then grbp<="111";
	end if;
	if (ll=103 and cc>=99 and cc<162) then grbp<="111";
	end if;
	if (ll=103 and cc>=186 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=103) then grbp<="111";
	end if;
	if (ll=103 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (ll=103 and cc>=237 and cc<240) then grbp<="111";
	end if;
	if (cc=61 and ll=104) then grbp<="111";
	end if;
	if (cc=98 and ll=104) then grbp<="111";
	end if;
	if (ll=104 and cc>=98 and cc<163) then grbp<="111";
	end if;
	if (ll=104 and cc>=185 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=104) then grbp<="111";
	end if;
	if (cc=190 and ll=104) then grbp<="111";
	end if;
	if (ll=104 and cc>=190 and cc<205) then grbp<="111";
	end if;
	if (cc=236 and ll=104) then grbp<="111";
	end if;
	if (ll=104 and cc>=236 and cc<238) then grbp<="111";
	end if;
	if (ll=105 and cc>=61 and cc<63) then grbp<="111";
	end if;
	if (ll=105 and cc>=98 and cc<163) then grbp<="111";
	end if;
	if (ll=105 and cc>=184 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=105) then grbp<="111";
	end if;
	if (ll=105 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=236 and ll=105) then grbp<="111";
	end if;
	if (ll=105 and cc>=236 and cc<238) then grbp<="111";
	end if;
	if (cc=97 and ll=106) then grbp<="111";
	end if;
	if (ll=106 and cc>=97 and cc<163) then grbp<="111";
	end if;
	if (ll=106 and cc>=184 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=106) then grbp<="111";
	end if;
	if (ll=106 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=236 and ll=106) then grbp<="111";
	end if;
	if (cc=238 and ll=106) then grbp<="111";
	end if;
	if (cc=243 and ll=106) then grbp<="111";
	end if;
	if (cc=245 and ll=106) then grbp<="111";
	end if;
	if (cc=61 and ll=107) then grbp<="111";
	end if;
	if (cc=96 and ll=107) then grbp<="111";
	end if;
	if (ll=107 and cc>=96 and cc<164) then grbp<="111";
	end if;
	if (ll=107 and cc>=183 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=107) then grbp<="111";
	end if;
	if (ll=107 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=235 and ll=107) then grbp<="111";
	end if;
	if (cc=249 and ll=107) then grbp<="111";
	end if;
	if (cc=61 and ll=108) then grbp<="111";
	end if;
	if (cc=97 and ll=108) then grbp<="111";
	end if;
	if (ll=108 and cc>=97 and cc<105) then grbp<="111";
	end if;
	if (ll=108 and cc>=107 and cc<165) then grbp<="111";
	end if;
	if (ll=108 and cc>=182 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=108) then grbp<="111";
	end if;
	if (ll=108 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=235 and ll=108) then grbp<="111";
	end if;
	if (cc=237 and ll=108) then grbp<="111";
	end if;
	if (ll=108 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (cc=60 and ll=109) then grbp<="111";
	end if;
	if (ll=109 and cc>=60 and cc<63) then grbp<="111";
	end if;
	if (cc=97 and ll=109) then grbp<="111";
	end if;
	if (ll=109 and cc>=97 and cc<99) then grbp<="111";
	end if;
	if (ll=109 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (ll=109 and cc>=106 and cc<166) then grbp<="111";
	end if;
	if (ll=109 and cc>=181 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=109) then grbp<="111";
	end if;
	if (ll=109 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=239 and ll=109) then grbp<="111";
	end if;
	if (cc=60 and ll=110) then grbp<="111";
	end if;
	if (ll=110 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=98 and ll=110) then grbp<="111";
	end if;
	if (cc=102 and ll=110) then grbp<="111";
	end if;
	if (ll=110 and cc>=102 and cc<104) then grbp<="111";
	end if;
	if (ll=110 and cc>=105 and cc<166) then grbp<="111";
	end if;
	if (ll=110 and cc>=180 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=110) then grbp<="111";
	end if;
	if (ll=110 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=234 and ll=110) then grbp<="111";
	end if;
	if (ll=110 and cc>=234 and cc<238) then grbp<="111";
	end if;
	if (ll=111 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (ll=111 and cc>=95 and cc<97) then grbp<="111";
	end if;
	if (cc=101 and ll=111) then grbp<="111";
	end if;
	if (ll=111 and cc>=101 and cc<103) then grbp<="111";
	end if;
	if (ll=111 and cc>=104 and cc<167) then grbp<="111";
	end if;
	if (ll=111 and cc>=179 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=111) then grbp<="111";
	end if;
	if (ll=111 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=234 and ll=111) then grbp<="111";
	end if;
	if (ll=111 and cc>=234 and cc<238) then grbp<="111";
	end if;
	if (cc=250 and ll=111) then grbp<="111";
	end if;
	if (cc=60 and ll=112) then grbp<="111";
	end if;
	if (ll=112 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=104 and ll=112) then grbp<="111";
	end if;
	if (ll=112 and cc>=104 and cc<167) then grbp<="111";
	end if;
	if (ll=112 and cc>=178 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=112) then grbp<="111";
	end if;
	if (ll=112 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (ll=112 and cc>=229 and cc<231) then grbp<="111";
	end if;
	if (cc=245 and ll=112) then grbp<="111";
	end if;
	if (cc=60 and ll=113) then grbp<="111";
	end if;
	if (ll=113 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (ll=113 and cc>=93 and cc<95) then grbp<="111";
	end if;
	if (cc=100 and ll=113) then grbp<="111";
	end if;
	if (cc=103 and ll=113) then grbp<="111";
	end if;
	if (ll=113 and cc>=103 and cc<167) then grbp<="111";
	end if;
	if (ll=113 and cc>=176 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=113) then grbp<="111";
	end if;
	if (ll=113 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=233 and ll=113) then grbp<="111";
	end if;
	if (cc=238 and ll=113) then grbp<="111";
	end if;
	if (ll=113 and cc>=238 and cc<240) then grbp<="111";
	end if;
	if (ll=114 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=103 and ll=114) then grbp<="111";
	end if;
	if (ll=114 and cc>=103 and cc<168) then grbp<="111";
	end if;
	if (ll=114 and cc>=175 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=114) then grbp<="111";
	end if;
	if (ll=114 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=240 and ll=114) then grbp<="111";
	end if;
	if (cc=60 and ll=115) then grbp<="111";
	end if;
	if (ll=115 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=98 and ll=115) then grbp<="111";
	end if;
	if (cc=102 and ll=115) then grbp<="111";
	end if;
	if (ll=115 and cc>=102 and cc<168) then grbp<="111";
	end if;
	if (ll=115 and cc>=174 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=115) then grbp<="111";
	end if;
	if (ll=115 and cc>=188 and cc<205) then grbp<="111";
	end if;
	if (cc=60 and ll=116) then grbp<="111";
	end if;
	if (ll=116 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=101 and ll=116) then grbp<="111";
	end if;
	if (ll=116 and cc>=101 and cc<104) then grbp<="111";
	end if;
	if (ll=116 and cc>=105 and cc<168) then grbp<="111";
	end if;
	if (ll=116 and cc>=173 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=116) then grbp<="111";
	end if;
	if (ll=116 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (cc=235 and ll=116) then grbp<="111";
	end if;
	if (cc=237 and ll=116) then grbp<="111";
	end if;
	if (cc=60 and ll=117) then grbp<="111";
	end if;
	if (cc=97 and ll=117) then grbp<="111";
	end if;
	if (cc=100 and ll=117) then grbp<="111";
	end if;
	if (ll=117 and cc>=100 and cc<118) then grbp<="111";
	end if;
	if (ll=117 and cc>=119 and cc<168) then grbp<="111";
	end if;
	if (ll=117 and cc>=172 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=117) then grbp<="111";
	end if;
	if (ll=117 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (cc=246 and ll=117) then grbp<="111";
	end if;
	if (cc=59 and ll=118) then grbp<="111";
	end if;
	if (ll=118 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=96 and ll=118) then grbp<="111";
	end if;
	if (cc=100 and ll=118) then grbp<="111";
	end if;
	if (cc=102 and ll=118) then grbp<="111";
	end if;
	if (ll=118 and cc>=102 and cc<169) then grbp<="111";
	end if;
	if (ll=118 and cc>=171 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=118) then grbp<="111";
	end if;
	if (ll=118 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (ll=118 and cc>=231 and cc<238) then grbp<="111";
	end if;
	if (cc=242 and ll=118) then grbp<="111";
	end if;
	if (cc=24 and ll=119) then grbp<="111";
	end if;
	if (cc=59 and ll=119) then grbp<="111";
	end if;
	if (ll=119 and cc>=59 and cc<62) then grbp<="111";
	end if;
	if (cc=100 and ll=119) then grbp<="111";
	end if;
	if (ll=119 and cc>=100 and cc<106) then grbp<="111";
	end if;
	if (ll=119 and cc>=107 and cc<169) then grbp<="111";
	end if;
	if (ll=119 and cc>=170 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=119) then grbp<="111";
	end if;
	if (ll=119 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (cc=235 and ll=119) then grbp<="111";
	end if;
	if (ll=119 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (cc=59 and ll=120) then grbp<="111";
	end if;
	if (ll=120 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=100 and ll=120) then grbp<="111";
	end if;
	if (ll=120 and cc>=100 and cc<115) then grbp<="111";
	end if;
	if (ll=120 and cc>=117 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=120) then grbp<="111";
	end if;
	if (ll=120 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (ll=120 and cc>=231 and cc<233) then grbp<="111";
	end if;
	if (ll=120 and cc>=236 and cc<238) then grbp<="111";
	end if;
	if (ll=121 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (ll=121 and cc>=101 and cc<115) then grbp<="111";
	end if;
	if (ll=121 and cc>=116 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=121) then grbp<="111";
	end if;
	if (ll=121 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (ll=121 and cc>=230 and cc<233) then grbp<="111";
	end if;
	if (ll=121 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (ll=122 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (ll=122 and cc>=101 and cc<103) then grbp<="111";
	end if;
	if (ll=122 and cc>=106 and cc<115) then grbp<="111";
	end if;
	if (ll=122 and cc>=116 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=122) then grbp<="111";
	end if;
	if (ll=122 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (ll=122 and cc>=229 and cc<231) then grbp<="111";
	end if;
	if (cc=236 and ll=122) then grbp<="111";
	end if;
	if (cc=238 and ll=122) then grbp<="111";
	end if;
	if (cc=59 and ll=123) then grbp<="111";
	end if;
	if (ll=123 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=102 and ll=123) then grbp<="111";
	end if;
	if (cc=105 and ll=123) then grbp<="111";
	end if;
	if (ll=123 and cc>=105 and cc<113) then grbp<="111";
	end if;
	if (ll=123 and cc>=115 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=123) then grbp<="111";
	end if;
	if (ll=123 and cc>=188 and cc<204) then grbp<="111";
	end if;
	if (ll=123 and cc>=229 and cc<237) then grbp<="111";
	end if;
	if (cc=241 and ll=123) then grbp<="111";
	end if;
	if (cc=245 and ll=123) then grbp<="111";
	end if;
	if (cc=59 and ll=124) then grbp<="111";
	end if;
	if (ll=124 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=103 and ll=124) then grbp<="111";
	end if;
	if (cc=105 and ll=124) then grbp<="111";
	end if;
	if (ll=124 and cc>=105 and cc<113) then grbp<="111";
	end if;
	if (ll=124 and cc>=114 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=124) then grbp<="111";
	end if;
	if (ll=124 and cc>=188 and cc<203) then grbp<="111";
	end if;
	if (ll=124 and cc>=230 and cc<232) then grbp<="111";
	end if;
	if (cc=238 and ll=124) then grbp<="111";
	end if;
	if (cc=241 and ll=124) then grbp<="111";
	end if;
	if (cc=243 and ll=124) then grbp<="111";
	end if;
	if (ll=124 and cc>=243 and cc<245) then grbp<="111";
	end if;
	if (cc=92 and ll=125) then grbp<="111";
	end if;
	if (cc=96 and ll=125) then grbp<="111";
	end if;
	if (cc=100 and ll=125) then grbp<="111";
	end if;
	if (cc=105 and ll=125) then grbp<="111";
	end if;
	if (ll=125 and cc>=105 and cc<111) then grbp<="111";
	end if;
	if (ll=125 and cc>=113 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=125) then grbp<="111";
	end if;
	if (ll=125 and cc>=188 and cc<203) then grbp<="111";
	end if;
	if (ll=125 and cc>=230 and cc<232) then grbp<="111";
	end if;
	if (cc=236 and ll=125) then grbp<="111";
	end if;
	if (cc=238 and ll=125) then grbp<="111";
	end if;
	if (cc=241 and ll=125) then grbp<="111";
	end if;
	if (ll=125 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (cc=59 and ll=126) then grbp<="111";
	end if;
	if (cc=62 and ll=126) then grbp<="111";
	end if;
	if (cc=91 and ll=126) then grbp<="111";
	end if;
	if (cc=99 and ll=126) then grbp<="111";
	end if;
	if (cc=104 and ll=126) then grbp<="111";
	end if;
	if (ll=126 and cc>=104 and cc<111) then grbp<="111";
	end if;
	if (ll=126 and cc>=112 and cc<117) then grbp<="111";
	end if;
	if (ll=126 and cc>=118 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=126) then grbp<="111";
	end if;
	if (ll=126 and cc>=188 and cc<203) then grbp<="111";
	end if;
	if (cc=228 and ll=126) then grbp<="111";
	end if;
	if (ll=126 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (ll=126 and cc>=232 and cc<236) then grbp<="111";
	end if;
	if (cc=59 and ll=127) then grbp<="111";
	end if;
	if (ll=127 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=107 and ll=127) then grbp<="111";
	end if;
	if (ll=127 and cc>=107 and cc<111) then grbp<="111";
	end if;
	if (ll=127 and cc>=112 and cc<118) then grbp<="111";
	end if;
	if (ll=127 and cc>=119 and cc<130) then grbp<="111";
	end if;
	if (ll=127 and cc>=131 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=127) then grbp<="111";
	end if;
	if (ll=127 and cc>=188 and cc<203) then grbp<="111";
	end if;
	if (ll=127 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=236 and ll=127) then grbp<="111";
	end if;
	if (cc=238 and ll=127) then grbp<="111";
	end if;
	if (cc=240 and ll=127) then grbp<="111";
	end if;
	if (cc=59 and ll=128) then grbp<="111";
	end if;
	if (cc=63 and ll=128) then grbp<="111";
	end if;
	if (cc=105 and ll=128) then grbp<="111";
	end if;
	if (ll=128 and cc>=105 and cc<109) then grbp<="111";
	end if;
	if (ll=128 and cc>=111 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=128) then grbp<="111";
	end if;
	if (ll=128 and cc>=188 and cc<203) then grbp<="111";
	end if;
	if (cc=227 and ll=128) then grbp<="111";
	end if;
	if (ll=128 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (ll=128 and cc>=231 and cc<233) then grbp<="111";
	end if;
	if (ll=128 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (cc=97 and ll=129) then grbp<="111";
	end if;
	if (cc=102 and ll=129) then grbp<="111";
	end if;
	if (ll=129 and cc>=102 and cc<104) then grbp<="111";
	end if;
	if (cc=108 and ll=129) then grbp<="111";
	end if;
	if (cc=110 and ll=129) then grbp<="111";
	end if;
	if (ll=129 and cc>=110 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=129) then grbp<="111";
	end if;
	if (ll=129 and cc>=188 and cc<202) then grbp<="111";
	end if;
	if (ll=129 and cc>=227 and cc<238) then grbp<="111";
	end if;
	if (ll=130 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=106 and ll=130) then grbp<="111";
	end if;
	if (ll=130 and cc>=106 and cc<108) then grbp<="111";
	end if;
	if (ll=130 and cc>=109 and cc<124) then grbp<="111";
	end if;
	if (ll=130 and cc>=125 and cc<132) then grbp<="111";
	end if;
	if (ll=130 and cc>=133 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=130) then grbp<="111";
	end if;
	if (ll=130 and cc>=188 and cc<197) then grbp<="111";
	end if;
	if (ll=130 and cc>=198 and cc<202) then grbp<="111";
	end if;
	if (ll=130 and cc>=227 and cc<231) then grbp<="111";
	end if;
	if (cc=234 and ll=130) then grbp<="111";
	end if;
	if (cc=236 and ll=130) then grbp<="111";
	end if;
	if (cc=249 and ll=130) then grbp<="111";
	end if;
	if (cc=59 and ll=131) then grbp<="111";
	end if;
	if (cc=61 and ll=131) then grbp<="111";
	end if;
	if (cc=88 and ll=131) then grbp<="111";
	end if;
	if (cc=95 and ll=131) then grbp<="111";
	end if;
	if (cc=100 and ll=131) then grbp<="111";
	end if;
	if (ll=131 and cc>=100 and cc<102) then grbp<="111";
	end if;
	if (ll=131 and cc>=109 and cc<132) then grbp<="111";
	end if;
	if (ll=131 and cc>=133 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=131) then grbp<="111";
	end if;
	if (ll=131 and cc>=188 and cc<192) then grbp<="111";
	end if;
	if (ll=131 and cc>=193 and cc<196) then grbp<="111";
	end if;
	if (ll=131 and cc>=198 and cc<202) then grbp<="111";
	end if;
	if (ll=131 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (cc=233 and ll=131) then grbp<="111";
	end if;
	if (ll=131 and cc>=233 and cc<236) then grbp<="111";
	end if;
	if (ll=131 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (cc=242 and ll=131) then grbp<="111";
	end if;
	if (cc=245 and ll=131) then grbp<="111";
	end if;
	if (cc=247 and ll=131) then grbp<="111";
	end if;
	if (cc=59 and ll=132) then grbp<="111";
	end if;
	if (cc=101 and ll=132) then grbp<="111";
	end if;
	if (cc=103 and ll=132) then grbp<="111";
	end if;
	if (cc=108 and ll=132) then grbp<="111";
	end if;
	if (cc=110 and ll=132) then grbp<="111";
	end if;
	if (ll=132 and cc>=110 and cc<122) then grbp<="111";
	end if;
	if (ll=132 and cc>=123 and cc<131) then grbp<="111";
	end if;
	if (ll=132 and cc>=132 and cc<155) then grbp<="111";
	end if;
	if (ll=132 and cc>=156 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=132) then grbp<="111";
	end if;
	if (ll=132 and cc>=188 and cc<196) then grbp<="111";
	end if;
	if (ll=132 and cc>=198 and cc<202) then grbp<="111";
	end if;
	if (ll=132 and cc>=226 and cc<237) then grbp<="111";
	end if;
	if (cc=250 and ll=132) then grbp<="111";
	end if;
	if (cc=59 and ll=133) then grbp<="111";
	end if;
	if (ll=133 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (ll=133 and cc>=103 and cc<105) then grbp<="111";
	end if;
	if (ll=133 and cc>=107 and cc<109) then grbp<="111";
	end if;
	if (ll=133 and cc>=110 and cc<130) then grbp<="111";
	end if;
	if (ll=133 and cc>=131 and cc<155) then grbp<="111";
	end if;
	if (ll=133 and cc>=156 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=133) then grbp<="111";
	end if;
	if (ll=133 and cc>=188 and cc<195) then grbp<="111";
	end if;
	if (ll=133 and cc>=197 and cc<201) then grbp<="111";
	end if;
	if (ll=133 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=133 and cc>=229 and cc<232) then grbp<="111";
	end if;
	if (cc=59 and ll=134) then grbp<="111";
	end if;
	if (cc=103 and ll=134) then grbp<="111";
	end if;
	if (ll=134 and cc>=103 and cc<105) then grbp<="111";
	end if;
	if (ll=134 and cc>=108 and cc<110) then grbp<="111";
	end if;
	if (ll=134 and cc>=111 and cc<123) then grbp<="111";
	end if;
	if (ll=134 and cc>=124 and cc<127) then grbp<="111";
	end if;
	if (ll=134 and cc>=129 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=134) then grbp<="111";
	end if;
	if (ll=134 and cc>=188 and cc<190) then grbp<="111";
	end if;
	if (ll=134 and cc>=191 and cc<194) then grbp<="111";
	end if;
	if (ll=134 and cc>=197 and cc<201) then grbp<="111";
	end if;
	if (ll=134 and cc>=225 and cc<232) then grbp<="111";
	end if;
	if (cc=237 and ll=134) then grbp<="111";
	end if;
	if (cc=58 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=106 and ll=135) then grbp<="111";
	end if;
	if (cc=109 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=109 and cc<111) then grbp<="111";
	end if;
	if (cc=115 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=115 and cc<117) then grbp<="111";
	end if;
	if (ll=135 and cc>=119 and cc<124) then grbp<="111";
	end if;
	if (cc=128 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=128 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=188 and cc<194) then grbp<="111";
	end if;
	if (ll=135 and cc>=196 and cc<201) then grbp<="111";
	end if;
	if (cc=226 and ll=135) then grbp<="111";
	end if;
	if (cc=228 and ll=135) then grbp<="111";
	end if;
	if (ll=135 and cc>=228 and cc<232) then grbp<="111";
	end if;
	if (cc=238 and ll=135) then grbp<="111";
	end if;
	if (cc=247 and ll=135) then grbp<="111";
	end if;
	if (cc=58 and ll=136) then grbp<="111";
	end if;
	if (cc=85 and ll=136) then grbp<="111";
	end if;
	if (cc=106 and ll=136) then grbp<="111";
	end if;
	if (ll=136 and cc>=106 and cc<108) then grbp<="111";
	end if;
	if (ll=136 and cc>=109 and cc<111) then grbp<="111";
	end if;
	if (ll=136 and cc>=113 and cc<117) then grbp<="111";
	end if;
	if (ll=136 and cc>=118 and cc<124) then grbp<="111";
	end if;
	if (ll=136 and cc>=128 and cc<140) then grbp<="111";
	end if;
	if (ll=136 and cc>=141 and cc<152) then grbp<="111";
	end if;
	if (ll=136 and cc>=153 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=136) then grbp<="111";
	end if;
	if (ll=136 and cc>=188 and cc<193) then grbp<="111";
	end if;
	if (ll=136 and cc>=195 and cc<201) then grbp<="111";
	end if;
	if (cc=225 and ll=136) then grbp<="111";
	end if;
	if (ll=136 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=235 and ll=136) then grbp<="111";
	end if;
	if (ll=136 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (cc=58 and ll=137) then grbp<="111";
	end if;
	if (cc=60 and ll=137) then grbp<="111";
	end if;
	if (cc=106 and ll=137) then grbp<="111";
	end if;
	if (ll=137 and cc>=106 and cc<108) then grbp<="111";
	end if;
	if (cc=114 and ll=137) then grbp<="111";
	end if;
	if (cc=116 and ll=137) then grbp<="111";
	end if;
	if (cc=118 and ll=137) then grbp<="111";
	end if;
	if (ll=137 and cc>=118 and cc<124) then grbp<="111";
	end if;
	if (ll=137 and cc>=126 and cc<150) then grbp<="111";
	end if;
	if (ll=137 and cc>=151 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=137) then grbp<="111";
	end if;
	if (ll=137 and cc>=188 and cc<193) then grbp<="111";
	end if;
	if (ll=137 and cc>=194 and cc<197) then grbp<="111";
	end if;
	if (ll=137 and cc>=198 and cc<201) then grbp<="111";
	end if;
	if (cc=225 and ll=137) then grbp<="111";
	end if;
	if (ll=137 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=137 and cc>=230 and cc<233) then grbp<="111";
	end if;
	if (cc=238 and ll=137) then grbp<="111";
	end if;
	if (cc=240 and ll=137) then grbp<="111";
	end if;
	if (cc=58 and ll=138) then grbp<="111";
	end if;
	if (ll=138 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=108 and ll=138) then grbp<="111";
	end if;
	if (cc=111 and ll=138) then grbp<="111";
	end if;
	if (ll=138 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (cc=118 and ll=138) then grbp<="111";
	end if;
	if (ll=138 and cc>=118 and cc<124) then grbp<="111";
	end if;
	if (ll=138 and cc>=125 and cc<150) then grbp<="111";
	end if;
	if (ll=138 and cc>=151 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=138) then grbp<="111";
	end if;
	if (ll=138 and cc>=188 and cc<192) then grbp<="111";
	end if;
	if (ll=138 and cc>=193 and cc<196) then grbp<="111";
	end if;
	if (ll=138 and cc>=198 and cc<200) then grbp<="111";
	end if;
	if (cc=224 and ll=138) then grbp<="111";
	end if;
	if (ll=138 and cc>=224 and cc<230) then grbp<="111";
	end if;
	if (cc=236 and ll=138) then grbp<="111";
	end if;
	if (cc=238 and ll=138) then grbp<="111";
	end if;
	if (cc=249 and ll=138) then grbp<="111";
	end if;
	if (cc=58 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=104 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=104 and cc<106) then grbp<="111";
	end if;
	if (cc=111 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (ll=139 and cc>=114 and cc<116) then grbp<="111";
	end if;
	if (cc=124 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=124 and cc<138) then grbp<="111";
	end if;
	if (ll=139 and cc>=139 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=188 and cc<191) then grbp<="111";
	end if;
	if (ll=139 and cc>=193 and cc<195) then grbp<="111";
	end if;
	if (ll=139 and cc>=197 and cc<200) then grbp<="111";
	end if;
	if (cc=236 and ll=139) then grbp<="111";
	end if;
	if (ll=139 and cc>=236 and cc<239) then grbp<="111";
	end if;
	if (cc=58 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=58 and cc<61) then grbp<="111";
	end if;
	if (cc=64 and ll=140) then grbp<="111";
	end if;
	if (cc=104 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=104 and cc<107) then grbp<="111";
	end if;
	if (cc=112 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=112 and cc<115) then grbp<="111";
	end if;
	if (cc=125 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=125 and cc<130) then grbp<="111";
	end if;
	if (ll=140 and cc>=131 and cc<145) then grbp<="111";
	end if;
	if (ll=140 and cc>=146 and cc<148) then grbp<="111";
	end if;
	if (ll=140 and cc>=149 and cc<188) then grbp<="111";
	end if;
	if (cc=189 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=189 and cc<191) then grbp<="111";
	end if;
	if (cc=197 and ll=140) then grbp<="111";
	end if;
	if (ll=140 and cc>=197 and cc<200) then grbp<="111";
	end if;
	if (cc=227 and ll=140) then grbp<="111";
	end if;
	if (cc=237 and ll=140) then grbp<="111";
	end if;
	if (cc=247 and ll=140) then grbp<="111";
	end if;
	if (cc=58 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=105 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=105 and cc<107) then grbp<="111";
	end if;
	if (cc=110 and ll=141) then grbp<="111";
	end if;
	if (cc=113 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=113 and cc<115) then grbp<="111";
	end if;
	if (ll=141 and cc>=123 and cc<125) then grbp<="111";
	end if;
	if (ll=141 and cc>=126 and cc<128) then grbp<="111";
	end if;
	if (ll=141 and cc>=130 and cc<137) then grbp<="111";
	end if;
	if (ll=141 and cc>=138 and cc<146) then grbp<="111";
	end if;
	if (cc=149 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=149 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=188 and cc<190) then grbp<="111";
	end if;
	if (cc=197 and ll=141) then grbp<="111";
	end if;
	if (ll=141 and cc>=197 and cc<200) then grbp<="111";
	end if;
	if (cc=225 and ll=141) then grbp<="111";
	end if;
	if (cc=232 and ll=141) then grbp<="111";
	end if;
	if (cc=248 and ll=141) then grbp<="111";
	end if;
	if (cc=58 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=65 and ll=142) then grbp<="111";
	end if;
	if (cc=106 and ll=142) then grbp<="111";
	end if;
	if (cc=115 and ll=142) then grbp<="111";
	end if;
	if (cc=118 and ll=142) then grbp<="111";
	end if;
	if (cc=123 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=123 and cc<129) then grbp<="111";
	end if;
	if (ll=142 and cc>=130 and cc<137) then grbp<="111";
	end if;
	if (cc=141 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=141 and cc<144) then grbp<="111";
	end if;
	if (cc=147 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=147 and cc<187) then grbp<="111";
	end if;
	if (cc=190 and ll=142) then grbp<="111";
	end if;
	if (cc=196 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=196 and cc<200) then grbp<="111";
	end if;
	if (cc=229 and ll=142) then grbp<="111";
	end if;
	if (ll=142 and cc>=229 and cc<232) then grbp<="111";
	end if;
	if (ll=142 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (cc=58 and ll=143) then grbp<="111";
	end if;
	if (ll=143 and cc>=58 and cc<61) then grbp<="111";
	end if;
	if (cc=120 and ll=143) then grbp<="111";
	end if;
	if (cc=125 and ll=143) then grbp<="111";
	end if;
	if (ll=143 and cc>=125 and cc<129) then grbp<="111";
	end if;
	if (ll=143 and cc>=134 and cc<137) then grbp<="111";
	end if;
	if (ll=143 and cc>=141 and cc<144) then grbp<="111";
	end if;
	if (cc=147 and ll=143) then grbp<="111";
	end if;
	if (ll=143 and cc>=147 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=143) then grbp<="111";
	end if;
	if (cc=196 and ll=143) then grbp<="111";
	end if;
	if (ll=143 and cc>=196 and cc<199) then grbp<="111";
	end if;
	if (ll=143 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (cc=235 and ll=143) then grbp<="111";
	end if;
	if (cc=58 and ll=144) then grbp<="111";
	end if;
	if (ll=144 and cc>=58 and cc<61) then grbp<="111";
	end if;
	if (cc=102 and ll=144) then grbp<="111";
	end if;
	if (cc=118 and ll=144) then grbp<="111";
	end if;
	if (ll=144 and cc>=118 and cc<121) then grbp<="111";
	end if;
	if (ll=144 and cc>=128 and cc<132) then grbp<="111";
	end if;
	if (cc=136 and ll=144) then grbp<="111";
	end if;
	if (ll=144 and cc>=136 and cc<138) then grbp<="111";
	end if;
	if (cc=146 and ll=144) then grbp<="111";
	end if;
	if (ll=144 and cc>=146 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=144) then grbp<="111";
	end if;
	if (cc=195 and ll=144) then grbp<="111";
	end if;
	if (ll=144 and cc>=195 and cc<199) then grbp<="111";
	end if;
	if (ll=144 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=232 and ll=144) then grbp<="111";
	end if;
	if (cc=240 and ll=144) then grbp<="111";
	end if;
	if (cc=245 and ll=144) then grbp<="111";
	end if;
	if (cc=58 and ll=145) then grbp<="111";
	end if;
	if (ll=145 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (ll=145 and cc>=61 and cc<63) then grbp<="111";
	end if;
	if (cc=118 and ll=145) then grbp<="111";
	end if;
	if (ll=145 and cc>=118 and cc<122) then grbp<="111";
	end if;
	if (ll=145 and cc>=129 and cc<133) then grbp<="111";
	end if;
	if (cc=143 and ll=145) then grbp<="111";
	end if;
	if (cc=146 and ll=145) then grbp<="111";
	end if;
	if (ll=145 and cc>=146 and cc<149) then grbp<="111";
	end if;
	if (ll=145 and cc>=150 and cc<188) then grbp<="111";
	end if;
	if (cc=195 and ll=145) then grbp<="111";
	end if;
	if (ll=145 and cc>=195 and cc<199) then grbp<="111";
	end if;
	if (cc=222 and ll=145) then grbp<="111";
	end if;
	if (ll=145 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=145 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=145 and cc>=233 and cc<235) then grbp<="111";
	end if;
	if (ll=145 and cc>=236 and cc<238) then grbp<="111";
	end if;
	if (ll=146 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=63 and ll=146) then grbp<="111";
	end if;
	if (cc=103 and ll=146) then grbp<="111";
	end if;
	if (cc=118 and ll=146) then grbp<="111";
	end if;
	if (ll=146 and cc>=118 and cc<122) then grbp<="111";
	end if;
	if (cc=143 and ll=146) then grbp<="111";
	end if;
	if (cc=145 and ll=146) then grbp<="111";
	end if;
	if (ll=146 and cc>=145 and cc<186) then grbp<="111";
	end if;
	if (ll=146 and cc>=195 and cc<198) then grbp<="111";
	end if;
	if (ll=146 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (cc=60 and ll=147) then grbp<="111";
	end if;
	if (cc=62 and ll=147) then grbp<="111";
	end if;
	if (cc=118 and ll=147) then grbp<="111";
	end if;
	if (ll=147 and cc>=118 and cc<121) then grbp<="111";
	end if;
	if (ll=147 and cc>=144 and cc<147) then grbp<="111";
	end if;
	if (ll=147 and cc>=148 and cc<185) then grbp<="111";
	end if;
	if (ll=147 and cc>=194 and cc<198) then grbp<="111";
	end if;
	if (cc=221 and ll=147) then grbp<="111";
	end if;
	if (ll=147 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=147 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (cc=233 and ll=147) then grbp<="111";
	end if;
	if (cc=237 and ll=147) then grbp<="111";
	end if;
	if (cc=239 and ll=147) then grbp<="111";
	end if;
	if (cc=58 and ll=148) then grbp<="111";
	end if;
	if (ll=148 and cc>=58 and cc<61) then grbp<="111";
	end if;
	if (cc=64 and ll=148) then grbp<="111";
	end if;
	if (cc=119 and ll=148) then grbp<="111";
	end if;
	if (ll=148 and cc>=119 and cc<121) then grbp<="111";
	end if;
	if (ll=148 and cc>=144 and cc<146) then grbp<="111";
	end if;
	if (ll=148 and cc>=148 and cc<184) then grbp<="111";
	end if;
	if (ll=148 and cc>=194 and cc<198) then grbp<="111";
	end if;
	if (ll=148 and cc>=221 and cc<228) then grbp<="111";
	end if;
	if (cc=233 and ll=148) then grbp<="111";
	end if;
	if (cc=235 and ll=148) then grbp<="111";
	end if;
	if (ll=148 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (ll=149 and cc>=58 and cc<60) then grbp<="111";
	end if;
	if (cc=63 and ll=149) then grbp<="111";
	end if;
	if (cc=119 and ll=149) then grbp<="111";
	end if;
	if (cc=143 and ll=149) then grbp<="111";
	end if;
	if (ll=149 and cc>=143 and cc<182) then grbp<="111";
	end if;
	if (ll=149 and cc>=193 and cc<197) then grbp<="111";
	end if;
	if (ll=149 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=149 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=231 and ll=149) then grbp<="111";
	end if;
	if (cc=233 and ll=149) then grbp<="111";
	end if;
	if (cc=235 and ll=149) then grbp<="111";
	end if;
	if (cc=59 and ll=150) then grbp<="111";
	end if;
	if (ll=150 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=143 and ll=150) then grbp<="111";
	end if;
	if (ll=150 and cc>=143 and cc<145) then grbp<="111";
	end if;
	if (ll=150 and cc>=146 and cc<181) then grbp<="111";
	end if;
	if (ll=150 and cc>=192 and cc<197) then grbp<="111";
	end if;
	if (ll=150 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (ll=150 and cc>=228 and cc<232) then grbp<="111";
	end if;
	if (ll=150 and cc>=233 and cc<236) then grbp<="111";
	end if;
	if (cc=59 and ll=151) then grbp<="111";
	end if;
	if (ll=151 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=64 and ll=151) then grbp<="111";
	end if;
	if (cc=142 and ll=151) then grbp<="111";
	end if;
	if (ll=151 and cc>=142 and cc<144) then grbp<="111";
	end if;
	if (ll=151 and cc>=145 and cc<179) then grbp<="111";
	end if;
	if (ll=151 and cc>=192 and cc<196) then grbp<="111";
	end if;
	if (ll=151 and cc>=220 and cc<224) then grbp<="111";
	end if;
	if (ll=151 and cc>=227 and cc<232) then grbp<="111";
	end if;
	if (ll=151 and cc>=233 and cc<236) then grbp<="111";
	end if;
	if (cc=245 and ll=151) then grbp<="111";
	end if;
	if (ll=151 and cc>=245 and cc<247) then grbp<="111";
	end if;
	if (ll=152 and cc>=59 and cc<63) then grbp<="111";
	end if;
	if (cc=141 and ll=152) then grbp<="111";
	end if;
	if (ll=152 and cc>=141 and cc<143) then grbp<="111";
	end if;
	if (ll=152 and cc>=145 and cc<178) then grbp<="111";
	end if;
	if (ll=152 and cc>=191 and cc<195) then grbp<="111";
	end if;
	if (ll=152 and cc>=220 and cc<223) then grbp<="111";
	end if;
	if (cc=227 and ll=152) then grbp<="111";
	end if;
	if (ll=152 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (ll=152 and cc>=232 and cc<239) then grbp<="111";
	end if;
	if (cc=244 and ll=152) then grbp<="111";
	end if;
	if (cc=59 and ll=153) then grbp<="111";
	end if;
	if (ll=153 and cc>=59 and cc<62) then grbp<="111";
	end if;
	if (cc=140 and ll=153) then grbp<="111";
	end if;
	if (ll=153 and cc>=140 and cc<142) then grbp<="111";
	end if;
	if (ll=153 and cc>=144 and cc<177) then grbp<="111";
	end if;
	if (ll=153 and cc>=190 and cc<194) then grbp<="111";
	end if;
	if (ll=153 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (cc=232 and ll=153) then grbp<="111";
	end if;
	if (ll=153 and cc>=232 and cc<234) then grbp<="111";
	end if;
	if (cc=237 and ll=153) then grbp<="111";
	end if;
	if (ll=153 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (cc=59 and ll=154) then grbp<="111";
	end if;
	if (ll=154 and cc>=59 and cc<65) then grbp<="111";
	end if;
	if (cc=143 and ll=154) then grbp<="111";
	end if;
	if (ll=154 and cc>=143 and cc<176) then grbp<="111";
	end if;
	if (ll=154 and cc>=189 and cc<194) then grbp<="111";
	end if;
	if (cc=221 and ll=154) then grbp<="111";
	end if;
	if (ll=154 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=154 and cc>=224 and cc<240) then grbp<="111";
	end if;
	if (ll=155 and cc>=59 and cc<61) then grbp<="111";
	end if;
	if (cc=64 and ll=155) then grbp<="111";
	end if;
	if (cc=139 and ll=155) then grbp<="111";
	end if;
	if (cc=143 and ll=155) then grbp<="111";
	end if;
	if (ll=155 and cc>=143 and cc<175) then grbp<="111";
	end if;
	if (ll=155 and cc>=188 and cc<193) then grbp<="111";
	end if;
	if (ll=155 and cc>=218 and cc<235) then grbp<="111";
	end if;
	if (cc=238 and ll=155) then grbp<="111";
	end if;
	if (cc=240 and ll=155) then grbp<="111";
	end if;
	if (cc=59 and ll=156) then grbp<="111";
	end if;
	if (cc=61 and ll=156) then grbp<="111";
	end if;
	if (ll=156 and cc>=61 and cc<64) then grbp<="111";
	end if;
	if (ll=156 and cc>=138 and cc<140) then grbp<="111";
	end if;
	if (ll=156 and cc>=142 and cc<174) then grbp<="111";
	end if;
	if (ll=156 and cc>=189 and cc<193) then grbp<="111";
	end if;
	if (ll=156 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=231 and ll=156) then grbp<="111";
	end if;
	if (cc=235 and ll=156) then grbp<="111";
	end if;
	if (ll=156 and cc>=235 and cc<239) then grbp<="111";
	end if;
	if (cc=249 and ll=156) then grbp<="111";
	end if;
	if (cc=59 and ll=157) then grbp<="111";
	end if;
	if (ll=157 and cc>=59 and cc<62) then grbp<="111";
	end if;
	if (cc=138 and ll=157) then grbp<="111";
	end if;
	if (cc=142 and ll=157) then grbp<="111";
	end if;
	if (ll=157 and cc>=142 and cc<173) then grbp<="111";
	end if;
	if (ll=157 and cc>=188 and cc<192) then grbp<="111";
	end if;
	if (ll=157 and cc>=219 and cc<237) then grbp<="111";
	end if;
	if (cc=245 and ll=157) then grbp<="111";
	end if;
	if (cc=248 and ll=157) then grbp<="111";
	end if;
	if (cc=60 and ll=158) then grbp<="111";
	end if;
	if (cc=62 and ll=158) then grbp<="111";
	end if;
	if (cc=64 and ll=158) then grbp<="111";
	end if;
	if (cc=137 and ll=158) then grbp<="111";
	end if;
	if (cc=141 and ll=158) then grbp<="111";
	end if;
	if (ll=158 and cc>=141 and cc<172) then grbp<="111";
	end if;
	if (ll=158 and cc>=188 and cc<192) then grbp<="111";
	end if;
	if (ll=158 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=232 and ll=158) then grbp<="111";
	end if;
	if (ll=158 and cc>=232 and cc<237) then grbp<="111";
	end if;
	if (cc=60 and ll=159) then grbp<="111";
	end if;
	if (ll=159 and cc>=60 and cc<63) then grbp<="111";
	end if;
	if (cc=136 and ll=159) then grbp<="111";
	end if;
	if (ll=159 and cc>=136 and cc<138) then grbp<="111";
	end if;
	if (ll=159 and cc>=140 and cc<171) then grbp<="111";
	end if;
	if (cc=188 and ll=159) then grbp<="111";
	end if;
	if (ll=159 and cc>=188 and cc<191) then grbp<="111";
	end if;
	if (cc=220 and ll=159) then grbp<="111";
	end if;
	if (ll=159 and cc>=220 and cc<239) then grbp<="111";
	end if;
	if (cc=242 and ll=159) then grbp<="111";
	end if;
	if (cc=60 and ll=160) then grbp<="111";
	end if;
	if (ll=160 and cc>=60 and cc<62) then grbp<="111";
	end if;
	if (cc=65 and ll=160) then grbp<="111";
	end if;
	if (cc=136 and ll=160) then grbp<="111";
	end if;
	if (cc=139 and ll=160) then grbp<="111";
	end if;
	if (ll=160 and cc>=139 and cc<170) then grbp<="111";
	end if;
	if (ll=160 and cc>=187 and cc<191) then grbp<="111";
	end if;
	if (cc=221 and ll=160) then grbp<="111";
	end if;
	if (cc=223 and ll=160) then grbp<="111";
	end if;
	if (ll=160 and cc>=223 and cc<235) then grbp<="111";
	end if;
	if (cc=240 and ll=160) then grbp<="111";
	end if;
	if (ll=160 and cc>=240 and cc<244) then grbp<="111";
	end if;
	if (cc=248 and ll=160) then grbp<="111";
	end if;
	if (cc=60 and ll=161) then grbp<="111";
	end if;
	if (ll=161 and cc>=60 and cc<65) then grbp<="111";
	end if;
	if (cc=139 and ll=161) then grbp<="111";
	end if;
	if (ll=161 and cc>=139 and cc<168) then grbp<="111";
	end if;
	if (cc=184 and ll=161) then grbp<="111";
	end if;
	if (ll=161 and cc>=184 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=161) then grbp<="111";
	end if;
	if (ll=161 and cc>=188 and cc<190) then grbp<="111";
	end if;
	if (ll=161 and cc>=218 and cc<230) then grbp<="111";
	end if;
	if (ll=161 and cc>=231 and cc<235) then grbp<="111";
	end if;
	if (ll=161 and cc>=236 and cc<240) then grbp<="111";
	end if;
	if (cc=244 and ll=161) then grbp<="111";
	end if;
	if (cc=60 and ll=162) then grbp<="111";
	end if;
	if (ll=162 and cc>=60 and cc<63) then grbp<="111";
	end if;
	if (cc=66 and ll=162) then grbp<="111";
	end if;
	if (cc=134 and ll=162) then grbp<="111";
	end if;
	if (ll=162 and cc>=134 and cc<136) then grbp<="111";
	end if;
	if (ll=162 and cc>=138 and cc<167) then grbp<="111";
	end if;
	if (cc=185 and ll=162) then grbp<="111";
	end if;
	if (ll=162 and cc>=185 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=162) then grbp<="111";
	end if;
	if (ll=162 and cc>=188 and cc<190) then grbp<="111";
	end if;
	if (ll=162 and cc>=217 and cc<239) then grbp<="111";
	end if;
	if (cc=243 and ll=162) then grbp<="111";
	end if;
	if (cc=247 and ll=162) then grbp<="111";
	end if;
	if (cc=61 and ll=163) then grbp<="111";
	end if;
	if (cc=63 and ll=163) then grbp<="111";
	end if;
	if (cc=65 and ll=163) then grbp<="111";
	end if;
	if (cc=137 and ll=163) then grbp<="111";
	end if;
	if (ll=163 and cc>=137 and cc<166) then grbp<="111";
	end if;
	if (cc=185 and ll=163) then grbp<="111";
	end if;
	if (ll=163 and cc>=185 and cc<188) then grbp<="111";
	end if;
	if (cc=188 and ll=163) then grbp<="111";
	end if;
	if (cc=217 and ll=163) then grbp<="111";
	end if;
	if (ll=163 and cc>=217 and cc<232) then grbp<="111";
	end if;
	if (ll=163 and cc>=234 and cc<236) then grbp<="111";
	end if;
	if (ll=163 and cc>=237 and cc<240) then grbp<="111";
	end if;
	if (ll=163 and cc>=241 and cc<244) then grbp<="111";
	end if;
	if (cc=61 and ll=164) then grbp<="111";
	end if;
	if (ll=164 and cc>=61 and cc<64) then grbp<="111";
	end if;
	if (cc=68 and ll=164) then grbp<="111";
	end if;
	if (cc=133 and ll=164) then grbp<="111";
	end if;
	if (cc=137 and ll=164) then grbp<="111";
	end if;
	if (ll=164 and cc>=137 and cc<165) then grbp<="111";
	end if;
	if (cc=184 and ll=164) then grbp<="111";
	end if;
	if (ll=164 and cc>=184 and cc<188) then grbp<="111";
	end if;
	if (cc=217 and ll=164) then grbp<="111";
	end if;
	if (cc=219 and ll=164) then grbp<="111";
	end if;
	if (ll=164 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (ll=164 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=164 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (ll=164 and cc>=232 and cc<239) then grbp<="111";
	end if;
	if (ll=164 and cc>=243 and cc<247) then grbp<="111";
	end if;
	if (ll=165 and cc>=61 and cc<65) then grbp<="111";
	end if;
	if (cc=131 and ll=165) then grbp<="111";
	end if;
	if (ll=165 and cc>=131 and cc<133) then grbp<="111";
	end if;
	if (ll=165 and cc>=136 and cc<165) then grbp<="111";
	end if;
	if (cc=177 and ll=165) then grbp<="111";
	end if;
	if (ll=165 and cc>=177 and cc<180) then grbp<="111";
	end if;
	if (cc=184 and ll=165) then grbp<="111";
	end if;
	if (ll=165 and cc>=184 and cc<188) then grbp<="111";
	end if;
	if (cc=217 and ll=165) then grbp<="111";
	end if;
	if (ll=165 and cc>=217 and cc<222) then grbp<="111";
	end if;
	if (ll=165 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=165 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=165 and cc>=231 and cc<234) then grbp<="111";
	end if;
	if (ll=165 and cc>=235 and cc<238) then grbp<="111";
	end if;
	if (ll=165 and cc>=239 and cc<241) then grbp<="111";
	end if;
	if (ll=165 and cc>=242 and cc<244) then grbp<="111";
	end if;
	if (ll=165 and cc>=246 and cc<248) then grbp<="111";
	end if;
	if (ll=166 and cc>=62 and cc<65) then grbp<="111";
	end if;
	if (ll=166 and cc>=131 and cc<133) then grbp<="111";
	end if;
	if (ll=166 and cc>=136 and cc<164) then grbp<="111";
	end if;
	if (ll=166 and cc>=183 and cc<187) then grbp<="111";
	end if;
	if (ll=166 and cc>=217 and cc<233) then grbp<="111";
	end if;
	if (ll=166 and cc>=235 and cc<239) then grbp<="111";
	end if;
	if (ll=166 and cc>=242 and cc<244) then grbp<="111";
	end if;
	if (cc=62 and ll=167) then grbp<="111";
	end if;
	if (ll=167 and cc>=62 and cc<64) then grbp<="111";
	end if;
	if (cc=69 and ll=167) then grbp<="111";
	end if;
	if (cc=127 and ll=167) then grbp<="111";
	end if;
	if (cc=131 and ll=167) then grbp<="111";
	end if;
	if (cc=135 and ll=167) then grbp<="111";
	end if;
	if (ll=167 and cc>=135 and cc<164) then grbp<="111";
	end if;
	if (ll=167 and cc>=182 and cc<186) then grbp<="111";
	end if;
	if (ll=167 and cc>=217 and cc<220) then grbp<="111";
	end if;
	if (cc=223 and ll=167) then grbp<="111";
	end if;
	if (ll=167 and cc>=223 and cc<230) then grbp<="111";
	end if;
	if (ll=167 and cc>=232 and cc<235) then grbp<="111";
	end if;
	if (ll=167 and cc>=236 and cc<243) then grbp<="111";
	end if;
	if (cc=246 and ll=167) then grbp<="111";
	end if;
	if (cc=250 and ll=167) then grbp<="111";
	end if;
	if (cc=62 and ll=168) then grbp<="111";
	end if;
	if (ll=168 and cc>=62 and cc<67) then grbp<="111";
	end if;
	if (cc=134 and ll=168) then grbp<="111";
	end if;
	if (ll=168 and cc>=134 and cc<164) then grbp<="111";
	end if;
	if (cc=181 and ll=168) then grbp<="111";
	end if;
	if (ll=168 and cc>=181 and cc<185) then grbp<="111";
	end if;
	if (ll=168 and cc>=216 and cc<221) then grbp<="111";
	end if;
	if (ll=168 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=168 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (ll=168 and cc>=231 and cc<239) then grbp<="111";
	end if;
	if (ll=168 and cc>=242 and cc<245) then grbp<="111";
	end if;
	if (cc=63 and ll=169) then grbp<="111";
	end if;
	if (ll=169 and cc>=63 and cc<67) then grbp<="111";
	end if;
	if (ll=169 and cc>=133 and cc<164) then grbp<="111";
	end if;
	if (ll=169 and cc>=180 and cc<184) then grbp<="111";
	end if;
	if (ll=169 and cc>=215 and cc<219) then grbp<="111";
	end if;
	if (ll=169 and cc>=220 and cc<224) then grbp<="111";
	end if;
	if (ll=169 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (ll=169 and cc>=231 and cc<239) then grbp<="111";
	end if;
	if (ll=169 and cc>=242 and cc<247) then grbp<="111";
	end if;
	if (ll=170 and cc>=63 and cc<68) then grbp<="111";
	end if;
	if (ll=170 and cc>=133 and cc<164) then grbp<="111";
	end if;
	if (ll=170 and cc>=179 and cc<184) then grbp<="111";
	end if;
	if (ll=170 and cc>=215 and cc<218) then grbp<="111";
	end if;
	if (ll=170 and cc>=220 and cc<223) then grbp<="111";
	end if;
	if (ll=170 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=170 and cc>=228 and cc<232) then grbp<="111";
	end if;
	if (ll=170 and cc>=233 and cc<240) then grbp<="111";
	end if;
	if (ll=170 and cc>=242 and cc<244) then grbp<="111";
	end if;
	if (ll=171 and cc>=63 and cc<68) then grbp<="111";
	end if;
	if (ll=171 and cc>=133 and cc<165) then grbp<="111";
	end if;
	if (ll=171 and cc>=178 and cc<183) then grbp<="111";
	end if;
	if (cc=217 and ll=171) then grbp<="111";
	end if;
	if (ll=171 and cc>=217 and cc<221) then grbp<="111";
	end if;
	if (ll=171 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=171 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=171 and cc>=230 and cc<237) then grbp<="111";
	end if;
	if (ll=171 and cc>=238 and cc<240) then grbp<="111";
	end if;
	if (ll=171 and cc>=242 and cc<244) then grbp<="111";
	end if;
	if (cc=249 and ll=171) then grbp<="111";
	end if;
	if (cc=64 and ll=172) then grbp<="111";
	end if;
	if (ll=172 and cc>=64 and cc<68) then grbp<="111";
	end if;
	if (cc=128 and ll=172) then grbp<="111";
	end if;
	if (cc=132 and ll=172) then grbp<="111";
	end if;
	if (ll=172 and cc>=132 and cc<165) then grbp<="111";
	end if;
	if (ll=172 and cc>=178 and cc<182) then grbp<="111";
	end if;
	if (ll=172 and cc>=214 and cc<236) then grbp<="111";
	end if;
	if (ll=172 and cc>=237 and cc<242) then grbp<="111";
	end if;
	if (cc=245 and ll=172) then grbp<="111";
	end if;
	if (cc=249 and ll=172) then grbp<="111";
	end if;
	if (cc=64 and ll=173) then grbp<="111";
	end if;
	if (ll=173 and cc>=64 and cc<68) then grbp<="111";
	end if;
	if (cc=131 and ll=173) then grbp<="111";
	end if;
	if (ll=173 and cc>=131 and cc<165) then grbp<="111";
	end if;
	if (ll=173 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=173 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (cc=223 and ll=173) then grbp<="111";
	end if;
	if (ll=173 and cc>=223 and cc<236) then grbp<="111";
	end if;
	if (cc=239 and ll=173) then grbp<="111";
	end if;
	if (ll=173 and cc>=239 and cc<242) then grbp<="111";
	end if;
	if (cc=247 and ll=173) then grbp<="111";
	end if;
	if (cc=64 and ll=174) then grbp<="111";
	end if;
	if (ll=174 and cc>=64 and cc<68) then grbp<="111";
	end if;
	if (cc=131 and ll=174) then grbp<="111";
	end if;
	if (ll=174 and cc>=131 and cc<165) then grbp<="111";
	end if;
	if (cc=214 and ll=174) then grbp<="111";
	end if;
	if (ll=174 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (ll=174 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=174 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (cc=233 and ll=174) then grbp<="111";
	end if;
	if (ll=174 and cc>=233 and cc<235) then grbp<="111";
	end if;
	if (ll=174 and cc>=237 and cc<241) then grbp<="111";
	end if;
	if (ll=174 and cc>=242 and cc<246) then grbp<="111";
	end if;
	if (cc=64 and ll=175) then grbp<="111";
	end if;
	if (ll=175 and cc>=64 and cc<70) then grbp<="111";
	end if;
	if (ll=175 and cc>=130 and cc<165) then grbp<="111";
	end if;
	if (cc=214 and ll=175) then grbp<="111";
	end if;
	if (ll=175 and cc>=214 and cc<224) then grbp<="111";
	end if;
	if (cc=227 and ll=175) then grbp<="111";
	end if;
	if (cc=229 and ll=175) then grbp<="111";
	end if;
	if (ll=175 and cc>=229 and cc<235) then grbp<="111";
	end if;
	if (ll=175 and cc>=236 and cc<241) then grbp<="111";
	end if;
	if (ll=175 and cc>=242 and cc<244) then grbp<="111";
	end if;
	if (cc=64 and ll=176) then grbp<="111";
	end if;
	if (ll=176 and cc>=64 and cc<69) then grbp<="111";
	end if;
	if (ll=176 and cc>=131 and cc<166) then grbp<="111";
	end if;
	if (cc=215 and ll=176) then grbp<="111";
	end if;
	if (ll=176 and cc>=215 and cc<218) then grbp<="111";
	end if;
	if (cc=221 and ll=176) then grbp<="111";
	end if;
	if (ll=176 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=176 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=176 and cc>=230 and cc<235) then grbp<="111";
	end if;
	if (ll=176 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (ll=176 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (ll=177 and cc>=64 and cc<70) then grbp<="111";
	end if;
	if (ll=177 and cc>=130 and cc<166) then grbp<="111";
	end if;
	if (cc=214 and ll=177) then grbp<="111";
	end if;
	if (ll=177 and cc>=214 and cc<220) then grbp<="111";
	end if;
	if (ll=177 and cc>=221 and cc<228) then grbp<="111";
	end if;
	if (ll=177 and cc>=229 and cc<238) then grbp<="111";
	end if;
	if (ll=177 and cc>=240 and cc<242) then grbp<="111";
	end if;
	if (cc=64 and ll=178) then grbp<="111";
	end if;
	if (ll=178 and cc>=64 and cc<69) then grbp<="111";
	end if;
	if (cc=130 and ll=178) then grbp<="111";
	end if;
	if (ll=178 and cc>=130 and cc<166) then grbp<="111";
	end if;
	if (cc=213 and ll=178) then grbp<="111";
	end if;
	if (ll=178 and cc>=213 and cc<222) then grbp<="111";
	end if;
	if (ll=178 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (ll=178 and cc>=229 and cc<238) then grbp<="111";
	end if;
	if (ll=179 and cc>=64 and cc<69) then grbp<="111";
	end if;
	if (ll=179 and cc>=128 and cc<166) then grbp<="111";
	end if;
	if (ll=179 and cc>=217 and cc<222) then grbp<="111";
	end if;
	if (cc=227 and ll=179) then grbp<="111";
	end if;
	if (cc=229 and ll=179) then grbp<="111";
	end if;
	if (ll=179 and cc>=229 and cc<233) then grbp<="111";
	end if;
	if (ll=179 and cc>=234 and cc<240) then grbp<="111";
	end if;
	if (ll=179 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (cc=247 and ll=179) then grbp<="111";
	end if;
	if (cc=64 and ll=180) then grbp<="111";
	end if;
	if (ll=180 and cc>=64 and cc<68) then grbp<="111";
	end if;
	if (ll=180 and cc>=128 and cc<166) then grbp<="111";
	end if;
	if (cc=215 and ll=180) then grbp<="111";
	end if;
	if (ll=180 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (ll=180 and cc>=218 and cc<222) then grbp<="111";
	end if;
	if (cc=227 and ll=180) then grbp<="111";
	end if;
	if (ll=180 and cc>=227 and cc<231) then grbp<="111";
	end if;
	if (ll=180 and cc>=234 and cc<236) then grbp<="111";
	end if;
	if (ll=180 and cc>=238 and cc<241) then grbp<="111";
	end if;
	if (cc=246 and ll=180) then grbp<="111";
	end if;
	if (cc=64 and ll=181) then grbp<="111";
	end if;
	if (ll=181 and cc>=64 and cc<69) then grbp<="111";
	end if;
	if (cc=128 and ll=181) then grbp<="111";
	end if;
	if (ll=181 and cc>=128 and cc<166) then grbp<="111";
	end if;
	if (ll=181 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=181 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=181) then grbp<="111";
	end if;
	if (ll=181 and cc>=218 and cc<224) then grbp<="111";
	end if;
	if (cc=227 and ll=181) then grbp<="111";
	end if;
	if (ll=181 and cc>=227 and cc<233) then grbp<="111";
	end if;
	if (ll=181 and cc>=234 and cc<239) then grbp<="111";
	end if;
	if (cc=242 and ll=181) then grbp<="111";
	end if;
	if (cc=244 and ll=181) then grbp<="111";
	end if;
	if (cc=246 and ll=181) then grbp<="111";
	end if;
	if (cc=64 and ll=182) then grbp<="111";
	end if;
	if (ll=182 and cc>=64 and cc<68) then grbp<="111";
	end if;
	if (cc=128 and ll=182) then grbp<="111";
	end if;
	if (ll=182 and cc>=128 and cc<166) then grbp<="111";
	end if;
	if (ll=182 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=182 and cc>=217 and cc<220) then grbp<="111";
	end if;
	if (ll=182 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=182 and cc>=229 and cc<231) then grbp<="111";
	end if;
	if (ll=182 and cc>=232 and cc<242) then grbp<="111";
	end if;
	if (cc=65 and ll=183) then grbp<="111";
	end if;
	if (ll=183 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (cc=125 and ll=183) then grbp<="111";
	end if;
	if (ll=183 and cc>=125 and cc<127) then grbp<="111";
	end if;
	if (ll=183 and cc>=129 and cc<167) then grbp<="111";
	end if;
	if (ll=183 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=183 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=183 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=183 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=183 and cc>=230 and cc<236) then grbp<="111";
	end if;
	if (ll=183 and cc>=237 and cc<240) then grbp<="111";
	end if;
	if (cc=65 and ll=184) then grbp<="111";
	end if;
	if (ll=184 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=184 and cc>=124 and cc<127) then grbp<="111";
	end if;
	if (ll=184 and cc>=129 and cc<167) then grbp<="111";
	end if;
	if (ll=184 and cc>=177 and cc<180) then grbp<="111";
	end if;
	if (cc=218 and ll=184) then grbp<="111";
	end if;
	if (cc=220 and ll=184) then grbp<="111";
	end if;
	if (ll=184 and cc>=220 and cc<225) then grbp<="111";
	end if;
	if (cc=229 and ll=184) then grbp<="111";
	end if;
	if (ll=184 and cc>=229 and cc<231) then grbp<="111";
	end if;
	if (ll=184 and cc>=234 and cc<236) then grbp<="111";
	end if;
	if (ll=184 and cc>=237 and cc<240) then grbp<="111";
	end if;
	if (cc=245 and ll=184) then grbp<="111";
	end if;
	if (cc=65 and ll=185) then grbp<="111";
	end if;
	if (ll=185 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (cc=124 and ll=185) then grbp<="111";
	end if;
	if (ll=185 and cc>=124 and cc<127) then grbp<="111";
	end if;
	if (ll=185 and cc>=129 and cc<143) then grbp<="111";
	end if;
	if (ll=185 and cc>=144 and cc<167) then grbp<="111";
	end if;
	if (ll=185 and cc>=177 and cc<180) then grbp<="111";
	end if;
	if (cc=216 and ll=185) then grbp<="111";
	end if;
	if (cc=218 and ll=185) then grbp<="111";
	end if;
	if (ll=185 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (cc=227 and ll=185) then grbp<="111";
	end if;
	if (ll=185 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=185 and cc>=233 and cc<239) then grbp<="111";
	end if;
	if (ll=185 and cc>=240 and cc<242) then grbp<="111";
	end if;
	if (cc=65 and ll=186) then grbp<="111";
	end if;
	if (ll=186 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=186 and cc>=123 and cc<128) then grbp<="111";
	end if;
	if (ll=186 and cc>=129 and cc<143) then grbp<="111";
	end if;
	if (ll=186 and cc>=144 and cc<167) then grbp<="111";
	end if;
	if (ll=186 and cc>=177 and cc<180) then grbp<="111";
	end if;
	if (cc=213 and ll=186) then grbp<="111";
	end if;
	if (ll=186 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=186) then grbp<="111";
	end if;
	if (ll=186 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (cc=226 and ll=186) then grbp<="111";
	end if;
	if (cc=228 and ll=186) then grbp<="111";
	end if;
	if (ll=186 and cc>=228 and cc<238) then grbp<="111";
	end if;
	if (cc=65 and ll=187) then grbp<="111";
	end if;
	if (ll=187 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=187 and cc>=123 and cc<128) then grbp<="111";
	end if;
	if (ll=187 and cc>=129 and cc<142) then grbp<="111";
	end if;
	if (ll=187 and cc>=144 and cc<167) then grbp<="111";
	end if;
	if (ll=187 and cc>=177 and cc<180) then grbp<="111";
	end if;
	if (cc=214 and ll=187) then grbp<="111";
	end if;
	if (cc=223 and ll=187) then grbp<="111";
	end if;
	if (ll=187 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=187 and cc>=229 and cc<233) then grbp<="111";
	end if;
	if (ll=187 and cc>=234 and cc<238) then grbp<="111";
	end if;
	if (cc=66 and ll=188) then grbp<="111";
	end if;
	if (ll=188 and cc>=66 and cc<68) then grbp<="111";
	end if;
	if (ll=188 and cc>=122 and cc<128) then grbp<="111";
	end if;
	if (ll=188 and cc>=129 and cc<141) then grbp<="111";
	end if;
	if (ll=188 and cc>=143 and cc<167) then grbp<="111";
	end if;
	if (ll=188 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=188 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (cc=228 and ll=188) then grbp<="111";
	end if;
	if (ll=188 and cc>=228 and cc<231) then grbp<="111";
	end if;
	if (ll=188 and cc>=232 and cc<240) then grbp<="111";
	end if;
	if (cc=247 and ll=188) then grbp<="111";
	end if;
	if (cc=249 and ll=188) then grbp<="111";
	end if;
	if (cc=66 and ll=189) then grbp<="111";
	end if;
	if (ll=189 and cc>=66 and cc<68) then grbp<="111";
	end if;
	if (ll=189 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=189 and cc>=129 and cc<141) then grbp<="111";
	end if;
	if (ll=189 and cc>=143 and cc<167) then grbp<="111";
	end if;
	if (ll=189 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=189 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (cc=216 and ll=189) then grbp<="111";
	end if;
	if (cc=232 and ll=189) then grbp<="111";
	end if;
	if (ll=189 and cc>=232 and cc<236) then grbp<="111";
	end if;
	if (cc=239 and ll=189) then grbp<="111";
	end if;
	if (ll=189 and cc>=239 and cc<241) then grbp<="111";
	end if;
	if (cc=249 and ll=189) then grbp<="111";
	end if;
	if (cc=66 and ll=190) then grbp<="111";
	end if;
	if (ll=190 and cc>=66 and cc<68) then grbp<="111";
	end if;
	if (ll=190 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=190 and cc>=129 and cc<140) then grbp<="111";
	end if;
	if (ll=190 and cc>=143 and cc<168) then grbp<="111";
	end if;
	if (ll=190 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=190 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (ll=190 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=190 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (cc=232 and ll=190) then grbp<="111";
	end if;
	if (ll=190 and cc>=232 and cc<237) then grbp<="111";
	end if;
	if (ll=190 and cc>=238 and cc<241) then grbp<="111";
	end if;
	if (ll=191 and cc>=66 and cc<68) then grbp<="111";
	end if;
	if (ll=191 and cc>=120 and cc<139) then grbp<="111";
	end if;
	if (ll=191 and cc>=142 and cc<168) then grbp<="111";
	end if;
	if (ll=191 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=191 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (cc=233 and ll=191) then grbp<="111";
	end if;
	if (ll=191 and cc>=233 and cc<236) then grbp<="111";
	end if;
	if (cc=241 and ll=191) then grbp<="111";
	end if;
	if (cc=67 and ll=192) then grbp<="111";
	end if;
	if (cc=120 and ll=192) then grbp<="111";
	end if;
	if (ll=192 and cc>=120 and cc<139) then grbp<="111";
	end if;
	if (ll=192 and cc>=141 and cc<168) then grbp<="111";
	end if;
	if (ll=192 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (cc=213 and ll=192) then grbp<="111";
	end if;
	if (cc=233 and ll=192) then grbp<="111";
	end if;
	if (cc=235 and ll=192) then grbp<="111";
	end if;
	if (cc=237 and ll=192) then grbp<="111";
	end if;
	if (ll=192 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (cc=242 and ll=192) then grbp<="111";
	end if;
	if (cc=246 and ll=192) then grbp<="111";
	end if;
	if (cc=67 and ll=193) then grbp<="111";
	end if;
	if (cc=119 and ll=193) then grbp<="111";
	end if;
	if (ll=193 and cc>=119 and cc<138) then grbp<="111";
	end if;
	if (ll=193 and cc>=141 and cc<168) then grbp<="111";
	end if;
	if (ll=193 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=193 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (cc=222 and ll=193) then grbp<="111";
	end if;
	if (cc=237 and ll=193) then grbp<="111";
	end if;
	if (ll=193 and cc>=237 and cc<239) then grbp<="111";
	end if;
	if (cc=67 and ll=194) then grbp<="111";
	end if;
	if (cc=112 and ll=194) then grbp<="111";
	end if;
	if (cc=119 and ll=194) then grbp<="111";
	end if;
	if (cc=121 and ll=194) then grbp<="111";
	end if;
	if (ll=194 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=194 and cc>=129 and cc<137) then grbp<="111";
	end if;
	if (ll=194 and cc>=140 and cc<168) then grbp<="111";
	end if;
	if (ll=194 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=194 and cc>=209 and cc<212) then grbp<="111";
	end if;
	if (cc=216 and ll=194) then grbp<="111";
	end if;
	if (cc=218 and ll=194) then grbp<="111";
	end if;
	if (ll=194 and cc>=218 and cc<224) then grbp<="111";
	end if;
	if (cc=238 and ll=194) then grbp<="111";
	end if;
	if (cc=22 and ll=195) then grbp<="111";
	end if;
	if (cc=118 and ll=195) then grbp<="111";
	end if;
	if (ll=195 and cc>=118 and cc<128) then grbp<="111";
	end if;
	if (ll=195 and cc>=129 and cc<137) then grbp<="111";
	end if;
	if (ll=195 and cc>=139 and cc<168) then grbp<="111";
	end if;
	if (ll=195 and cc>=178 and cc<180) then grbp<="111";
	end if;
	if (ll=195 and cc>=209 and cc<213) then grbp<="111";
	end if;
	if (cc=216 and ll=195) then grbp<="111";
	end if;
	if (cc=218 and ll=195) then grbp<="111";
	end if;
	if (ll=195 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (cc=224 and ll=195) then grbp<="111";
	end if;
	if (cc=241 and ll=195) then grbp<="111";
	end if;
	if (ll=195 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (cc=118 and ll=196) then grbp<="111";
	end if;
	if (cc=121 and ll=196) then grbp<="111";
	end if;
	if (ll=196 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=196 and cc>=129 and cc<136) then grbp<="111";
	end if;
	if (cc=139 and ll=196) then grbp<="111";
	end if;
	if (ll=196 and cc>=139 and cc<168) then grbp<="111";
	end if;
	if (cc=209 and ll=196) then grbp<="111";
	end if;
	if (cc=211 and ll=196) then grbp<="111";
	end if;
	if (ll=196 and cc>=211 and cc<217) then grbp<="111";
	end if;
	if (ll=196 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=196 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (cc=233 and ll=196) then grbp<="111";
	end if;
	if (cc=117 and ll=197) then grbp<="111";
	end if;
	if (ll=197 and cc>=117 and cc<119) then grbp<="111";
	end if;
	if (ll=197 and cc>=121 and cc<135) then grbp<="111";
	end if;
	if (ll=197 and cc>=136 and cc<169) then grbp<="111";
	end if;
	if (cc=209 and ll=197) then grbp<="111";
	end if;
	if (cc=211 and ll=197) then grbp<="111";
	end if;
	if (cc=213 and ll=197) then grbp<="111";
	end if;
	if (ll=197 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=197 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=197 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (cc=244 and ll=197) then grbp<="111";
	end if;
	if (cc=117 and ll=198) then grbp<="111";
	end if;
	if (cc=120 and ll=198) then grbp<="111";
	end if;
	if (ll=198 and cc>=120 and cc<134) then grbp<="111";
	end if;
	if (ll=198 and cc>=135 and cc<169) then grbp<="111";
	end if;
	if (cc=209 and ll=198) then grbp<="111";
	end if;
	if (ll=198 and cc>=209 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=198) then grbp<="111";
	end if;
	if (ll=198 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (cc=229 and ll=198) then grbp<="111";
	end if;
	if (cc=232 and ll=198) then grbp<="111";
	end if;
	if (cc=244 and ll=198) then grbp<="111";
	end if;
	if (cc=116 and ll=199) then grbp<="111";
	end if;
	if (ll=199 and cc>=116 and cc<120) then grbp<="111";
	end if;
	if (ll=199 and cc>=121 and cc<133) then grbp<="111";
	end if;
	if (ll=199 and cc>=134 and cc<169) then grbp<="111";
	end if;
	if (ll=199 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (ll=199 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (cc=219 and ll=199) then grbp<="111";
	end if;
	if (ll=199 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=23 and ll=200) then grbp<="111";
	end if;
	if (cc=69 and ll=200) then grbp<="111";
	end if;
	if (cc=116 and ll=200) then grbp<="111";
	end if;
	if (cc=118 and ll=200) then grbp<="111";
	end if;
	if (ll=200 and cc>=118 and cc<132) then grbp<="111";
	end if;
	if (ll=200 and cc>=134 and cc<169) then grbp<="111";
	end if;
	if (ll=200 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=212 and ll=200) then grbp<="111";
	end if;
	if (ll=200 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=219 and ll=200) then grbp<="111";
	end if;
	if (ll=200 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=201 and cc>=115 and cc<131) then grbp<="111";
	end if;
	if (ll=201 and cc>=136 and cc<169) then grbp<="111";
	end if;
	if (ll=201 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=210 and ll=201) then grbp<="111";
	end if;
	if (ll=201 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=201 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (cc=63 and ll=202) then grbp<="111";
	end if;
	if (cc=115 and ll=202) then grbp<="111";
	end if;
	if (ll=202 and cc>=115 and cc<121) then grbp<="111";
	end if;
	if (ll=202 and cc>=122 and cc<130) then grbp<="111";
	end if;
	if (ll=202 and cc>=137 and cc<169) then grbp<="111";
	end if;
	if (ll=202 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=211 and ll=202) then grbp<="111";
	end if;
	if (cc=213 and ll=202) then grbp<="111";
	end if;
	if (ll=202 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=202 and cc>=220 and cc<225) then grbp<="111";
	end if;
	if (cc=62 and ll=203) then grbp<="111";
	end if;
	if (cc=115 and ll=203) then grbp<="111";
	end if;
	if (ll=203 and cc>=115 and cc<129) then grbp<="111";
	end if;
	if (ll=203 and cc>=139 and cc<168) then grbp<="111";
	end if;
	if (ll=203 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (ll=203 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (ll=203 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (cc=234 and ll=203) then grbp<="111";
	end if;
	if (cc=236 and ll=203) then grbp<="111";
	end if;
	if (cc=239 and ll=203) then grbp<="111";
	end if;
	if (cc=62 and ll=204) then grbp<="111";
	end if;
	if (cc=71 and ll=204) then grbp<="111";
	end if;
	if (cc=114 and ll=204) then grbp<="111";
	end if;
	if (cc=116 and ll=204) then grbp<="111";
	end if;
	if (ll=204 and cc>=116 and cc<120) then grbp<="111";
	end if;
	if (ll=204 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=204 and cc>=140 and cc<168) then grbp<="111";
	end if;
	if (ll=204 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=210 and ll=204) then grbp<="111";
	end if;
	if (cc=214 and ll=204) then grbp<="111";
	end if;
	if (cc=222 and ll=204) then grbp<="111";
	end if;
	if (cc=231 and ll=204) then grbp<="111";
	end if;
	if (cc=237 and ll=204) then grbp<="111";
	end if;
	if (cc=239 and ll=204) then grbp<="111";
	end if;
	if (cc=62 and ll=205) then grbp<="111";
	end if;
	if (cc=70 and ll=205) then grbp<="111";
	end if;
	if (ll=205 and cc>=70 and cc<73) then grbp<="111";
	end if;
	if (ll=205 and cc>=114 and cc<120) then grbp<="111";
	end if;
	if (ll=205 and cc>=121 and cc<128) then grbp<="111";
	end if;
	if (ll=205 and cc>=141 and cc<167) then grbp<="111";
	end if;
	if (ll=205 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=217 and ll=205) then grbp<="111";
	end if;
	if (cc=221 and ll=205) then grbp<="111";
	end if;
	if (ll=205 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (cc=236 and ll=205) then grbp<="111";
	end if;
	if (ll=205 and cc>=236 and cc<240) then grbp<="111";
	end if;
	if (cc=62 and ll=206) then grbp<="111";
	end if;
	if (cc=70 and ll=206) then grbp<="111";
	end if;
	if (cc=113 and ll=206) then grbp<="111";
	end if;
	if (cc=115 and ll=206) then grbp<="111";
	end if;
	if (ll=206 and cc>=115 and cc<127) then grbp<="111";
	end if;
	if (ll=206 and cc>=142 and cc<166) then grbp<="111";
	end if;
	if (ll=206 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=219 and ll=206) then grbp<="111";
	end if;
	if (cc=221 and ll=206) then grbp<="111";
	end if;
	if (ll=206 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (ll=206 and cc>=235 and cc<239) then grbp<="111";
	end if;
	if (cc=70 and ll=207) then grbp<="111";
	end if;
	if (cc=113 and ll=207) then grbp<="111";
	end if;
	if (cc=115 and ll=207) then grbp<="111";
	end if;
	if (ll=207 and cc>=115 and cc<126) then grbp<="111";
	end if;
	if (ll=207 and cc>=143 and cc<163) then grbp<="111";
	end if;
	if (ll=207 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (ll=207 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=226 and ll=207) then grbp<="111";
	end if;
	if (cc=234 and ll=207) then grbp<="111";
	end if;
	if (ll=207 and cc>=234 and cc<239) then grbp<="111";
	end if;
	if (cc=112 and ll=208) then grbp<="111";
	end if;
	if (ll=208 and cc>=112 and cc<114) then grbp<="111";
	end if;
	if (ll=208 and cc>=115 and cc<125) then grbp<="111";
	end if;
	if (cc=145 and ll=208) then grbp<="111";
	end if;
	if (ll=208 and cc>=145 and cc<162) then grbp<="111";
	end if;
	if (ll=208 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=215 and ll=208) then grbp<="111";
	end if;
	if (cc=217 and ll=208) then grbp<="111";
	end if;
	if (cc=220 and ll=208) then grbp<="111";
	end if;
	if (cc=223 and ll=208) then grbp<="111";
	end if;
	if (cc=231 and ll=208) then grbp<="111";
	end if;
	if (cc=234 and ll=208) then grbp<="111";
	end if;
	if (ll=208 and cc>=234 and cc<239) then grbp<="111";
	end if;
	if (ll=208 and cc>=240 and cc<242) then grbp<="111";
	end if;
	if (cc=114 and ll=209) then grbp<="111";
	end if;
	if (ll=209 and cc>=114 and cc<119) then grbp<="111";
	end if;
	if (ll=209 and cc>=120 and cc<125) then grbp<="111";
	end if;
	if (cc=145 and ll=209) then grbp<="111";
	end if;
	if (ll=209 and cc>=145 and cc<161) then grbp<="111";
	end if;
	if (ll=209 and cc>=179 and cc<181) then grbp<="111";
	end if;
	if (cc=211 and ll=209) then grbp<="111";
	end if;
	if (cc=213 and ll=209) then grbp<="111";
	end if;
	if (cc=223 and ll=209) then grbp<="111";
	end if;
	if (cc=235 and ll=209) then grbp<="111";
	end if;
	if (cc=237 and ll=209) then grbp<="111";
	end if;
	if (ll=209 and cc>=237 and cc<242) then grbp<="111";
	end if;
	if (ll=210 and cc>=111 and cc<124) then grbp<="111";
	end if;
	if (ll=210 and cc>=146 and cc<161) then grbp<="111";
	end if;
	if (cc=234 and ll=210) then grbp<="111";
	end if;
	if (cc=237 and ll=210) then grbp<="111";
	end if;
	if (ll=210 and cc>=237 and cc<242) then grbp<="111";
	end if;
	if (ll=210 and cc>=243 and cc<245) then grbp<="111";
	end if;
	if (cc=111 and ll=211) then grbp<="111";
	end if;
	if (ll=211 and cc>=111 and cc<113) then grbp<="111";
	end if;
	if (ll=211 and cc>=114 and cc<123) then grbp<="111";
	end if;
	if (ll=211 and cc>=148 and cc<160) then grbp<="111";
	end if;
	if (cc=209 and ll=211) then grbp<="111";
	end if;
	if (cc=234 and ll=211) then grbp<="111";
	end if;
	if (cc=237 and ll=211) then grbp<="111";
	end if;
	if (ll=211 and cc>=237 and cc<242) then grbp<="111";
	end if;
	if (ll=211 and cc>=243 and cc<245) then grbp<="111";
	end if;
	if (cc=110 and ll=212) then grbp<="111";
	end if;
	if (ll=212 and cc>=110 and cc<123) then grbp<="111";
	end if;
	if (cc=150 and ll=212) then grbp<="111";
	end if;
	if (ll=212 and cc>=150 and cc<160) then grbp<="111";
	end if;
	if (cc=221 and ll=212) then grbp<="111";
	end if;
	if (cc=238 and ll=212) then grbp<="111";
	end if;
	if (ll=212 and cc>=238 and cc<240) then grbp<="111";
	end if;
	if (ll=212 and cc>=243 and cc<246) then grbp<="111";
	end if;
	if (cc=110 and ll=213) then grbp<="111";
	end if;
	if (ll=213 and cc>=110 and cc<122) then grbp<="111";
	end if;
	if (ll=213 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (cc=206 and ll=213) then grbp<="111";
	end if;
	if (cc=208 and ll=213) then grbp<="111";
	end if;
	if (cc=231 and ll=213) then grbp<="111";
	end if;
	if (cc=236 and ll=213) then grbp<="111";
	end if;
	if (ll=213 and cc>=236 and cc<240) then grbp<="111";
	end if;
	if (ll=213 and cc>=243 and cc<245) then grbp<="111";
	end if;
	if (cc=110 and ll=214) then grbp<="111";
	end if;
	if (ll=214 and cc>=110 and cc<121) then grbp<="111";
	end if;
	if (ll=214 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (cc=209 and ll=214) then grbp<="111";
	end if;
	if (cc=235 and ll=214) then grbp<="111";
	end if;
	if (cc=237 and ll=214) then grbp<="111";
	end if;
	if (cc=239 and ll=214) then grbp<="111";
	end if;
	if (ll=214 and cc>=239 and cc<241) then grbp<="111";
	end if;
	if (ll=215 and cc>=54 and cc<56) then grbp<="111";
	end if;
	if (ll=215 and cc>=109 and cc<121) then grbp<="111";
	end if;
	if (ll=215 and cc>=150 and cc<158) then grbp<="111";
	end if;
	if (cc=208 and ll=215) then grbp<="111";
	end if;
	if (cc=213 and ll=215) then grbp<="111";
	end if;
	if (cc=234 and ll=215) then grbp<="111";
	end if;
	if (cc=236 and ll=215) then grbp<="111";
	end if;
	if (cc=54 and ll=216) then grbp<="111";
	end if;
	if (ll=216 and cc>=54 and cc<56) then grbp<="111";
	end if;
	if (cc=111 and ll=216) then grbp<="111";
	end if;
	if (ll=216 and cc>=111 and cc<120) then grbp<="111";
	end if;
	if (ll=216 and cc>=150 and cc<158) then grbp<="111";
	end if;
	if (cc=233 and ll=216) then grbp<="111";
	end if;
	if (ll=216 and cc>=233 and cc<235) then grbp<="111";
	end if;
	if (cc=53 and ll=217) then grbp<="111";
	end if;
	if (ll=217 and cc>=53 and cc<55) then grbp<="111";
	end if;
	if (ll=217 and cc>=108 and cc<120) then grbp<="111";
	end if;
	if (ll=217 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (cc=204 and ll=217) then grbp<="111";
	end if;
	if (cc=235 and ll=217) then grbp<="111";
	end if;
	if (ll=217 and cc>=235 and cc<237) then grbp<="111";
	end if;
	if (cc=52 and ll=218) then grbp<="111";
	end if;
	if (ll=218 and cc>=52 and cc<55) then grbp<="111";
	end if;
	if (cc=108 and ll=218) then grbp<="111";
	end if;
	if (ll=218 and cc>=108 and cc<119) then grbp<="111";
	end if;
	if (ll=218 and cc>=133 and cc<135) then grbp<="111";
	end if;
	if (ll=218 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (cc=180 and ll=218) then grbp<="111";
	end if;
	if (ll=218 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=237 and ll=218) then grbp<="111";
	end if;
	if (cc=52 and ll=219) then grbp<="111";
	end if;
	if (ll=219 and cc>=52 and cc<55) then grbp<="111";
	end if;
	if (ll=219 and cc>=108 and cc<118) then grbp<="111";
	end if;
	if (ll=219 and cc>=133 and cc<137) then grbp<="111";
	end if;
	if (ll=219 and cc>=150 and cc<156) then grbp<="111";
	end if;
	if (cc=180 and ll=219) then grbp<="111";
	end if;
	if (ll=219 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=236 and ll=219) then grbp<="111";
	end if;
	if (cc=238 and ll=219) then grbp<="111";
	end if;
	if (cc=24 and ll=220) then grbp<="111";
	end if;
	if (cc=53 and ll=220) then grbp<="111";
	end if;
	if (ll=220 and cc>=53 and cc<55) then grbp<="111";
	end if;
	if (ll=220 and cc>=107 and cc<118) then grbp<="111";
	end if;
	if (ll=220 and cc>=133 and cc<137) then grbp<="111";
	end if;
	if (ll=220 and cc>=150 and cc<156) then grbp<="111";
	end if;
	if (ll=220 and cc>=164 and cc<166) then grbp<="111";
	end if;
	if (cc=237 and ll=220) then grbp<="111";
	end if;
	if (cc=26 and ll=221) then grbp<="111";
	end if;
	if (cc=53 and ll=221) then grbp<="111";
	end if;
	if (ll=221 and cc>=53 and cc<56) then grbp<="111";
	end if;
	if (ll=221 and cc>=107 and cc<118) then grbp<="111";
	end if;
	if (ll=221 and cc>=133 and cc<138) then grbp<="111";
	end if;
	if (ll=221 and cc>=150 and cc<155) then grbp<="111";
	end if;
	if (cc=180 and ll=221) then grbp<="111";
	end if;
	if (ll=221 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=56 and ll=222) then grbp<="111";
	end if;
	if (ll=222 and cc>=56 and cc<58) then grbp<="111";
	end if;
	if (ll=222 and cc>=107 and cc<117) then grbp<="111";
	end if;
	if (ll=222 and cc>=133 and cc<138) then grbp<="111";
	end if;
	if (ll=222 and cc>=150 and cc<155) then grbp<="111";
	end if;
	if (ll=222 and cc>=164 and cc<166) then grbp<="111";
	end if;
	if (ll=222 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=208 and ll=222) then grbp<="111";
	end if;
	if (cc=25 and ll=223) then grbp<="111";
	end if;
	if (cc=53 and ll=223) then grbp<="111";
	end if;
	if (cc=56 and ll=223) then grbp<="111";
	end if;
	if (ll=223 and cc>=56 and cc<58) then grbp<="111";
	end if;
	if (ll=223 and cc>=107 and cc<116) then grbp<="111";
	end if;
	if (ll=223 and cc>=133 and cc<138) then grbp<="111";
	end if;
	if (ll=223 and cc>=149 and cc<155) then grbp<="111";
	end if;
	if (ll=223 and cc>=164 and cc<166) then grbp<="111";
	end if;
	if (ll=223 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=249 and ll=223) then grbp<="111";
	end if;
	if (ll=223 and cc>=249 and cc<251) then grbp<="111";
	end if;
	if (cc=56 and ll=224) then grbp<="111";
	end if;
	if (ll=224 and cc>=56 and cc<59) then grbp<="111";
	end if;
	if (ll=224 and cc>=106 and cc<116) then grbp<="111";
	end if;
	if (ll=224 and cc>=132 and cc<138) then grbp<="111";
	end if;
	if (ll=224 and cc>=149 and cc<155) then grbp<="111";
	end if;
	if (ll=224 and cc>=164 and cc<166) then grbp<="111";
	end if;
	if (ll=224 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=248 and ll=224) then grbp<="111";
	end if;
	if (ll=224 and cc>=248 and cc<251) then grbp<="111";
	end if;
	if (cc=53 and ll=225) then grbp<="111";
	end if;
	if (cc=55 and ll=225) then grbp<="111";
	end if;
	if (ll=225 and cc>=55 and cc<60) then grbp<="111";
	end if;
	if (cc=108 and ll=225) then grbp<="111";
	end if;
	if (ll=225 and cc>=108 and cc<115) then grbp<="111";
	end if;
	if (ll=225 and cc>=132 and cc<137) then grbp<="111";
	end if;
	if (ll=225 and cc>=150 and cc<155) then grbp<="111";
	end if;
	if (ll=225 and cc>=163 and cc<166) then grbp<="111";
	end if;
	if (ll=225 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=248 and ll=225) then grbp<="111";
	end if;
	if (ll=225 and cc>=248 and cc<251) then grbp<="111";
	end if;
	if (cc=53 and ll=226) then grbp<="111";
	end if;
	if (cc=55 and ll=226) then grbp<="111";
	end if;
	if (ll=226 and cc>=55 and cc<59) then grbp<="111";
	end if;
	if (ll=226 and cc>=105 and cc<107) then grbp<="111";
	end if;
	if (ll=226 and cc>=108 and cc<115) then grbp<="111";
	end if;
	if (ll=226 and cc>=131 and cc<137) then grbp<="111";
	end if;
	if (ll=226 and cc>=150 and cc<155) then grbp<="111";
	end if;
	if (ll=226 and cc>=163 and cc<166) then grbp<="111";
	end if;
	if (ll=226 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=246 and ll=226) then grbp<="111";
	end if;
	if (ll=226 and cc>=246 and cc<251) then grbp<="111";
	end if;
	if (cc=53 and ll=227) then grbp<="111";
	end if;
	if (ll=227 and cc>=53 and cc<58) then grbp<="111";
	end if;
	if (ll=227 and cc>=105 and cc<114) then grbp<="111";
	end if;
	if (ll=227 and cc>=131 and cc<137) then grbp<="111";
	end if;
	if (ll=227 and cc>=149 and cc<155) then grbp<="111";
	end if;
	if (ll=227 and cc>=162 and cc<165) then grbp<="111";
	end if;
	if (ll=227 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (ll=227 and cc>=202 and cc<204) then grbp<="111";
	end if;
	if (ll=227 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=246 and ll=227) then grbp<="111";
	end if;
	if (ll=227 and cc>=246 and cc<251) then grbp<="111";
	end if;
	if (cc=25 and ll=228) then grbp<="111";
	end if;
	if (cc=51 and ll=228) then grbp<="111";
	end if;
	if (cc=53 and ll=228) then grbp<="111";
	end if;
	if (ll=228 and cc>=53 and cc<57) then grbp<="111";
	end if;
	if (ll=228 and cc>=105 and cc<113) then grbp<="111";
	end if;
	if (ll=228 and cc>=131 and cc<138) then grbp<="111";
	end if;
	if (ll=228 and cc>=150 and cc<155) then grbp<="111";
	end if;
	if (ll=228 and cc>=162 and cc<164) then grbp<="111";
	end if;
	if (ll=228 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (ll=228 and cc>=202 and cc<204) then grbp<="111";
	end if;
	if (ll=228 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=228 and cc>=245 and cc<251) then grbp<="111";
	end if;
	if (cc=50 and ll=229) then grbp<="111";
	end if;
	if (cc=52 and ll=229) then grbp<="111";
	end if;
	if (cc=54 and ll=229) then grbp<="111";
	end if;
	if (ll=229 and cc>=54 and cc<56) then grbp<="111";
	end if;
	if (ll=229 and cc>=104 and cc<113) then grbp<="111";
	end if;
	if (ll=229 and cc>=134 and cc<140) then grbp<="111";
	end if;
	if (ll=229 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (ll=229 and cc>=162 and cc<164) then grbp<="111";
	end if;
	if (ll=229 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=213 and ll=229) then grbp<="111";
	end if;
	if (cc=216 and ll=229) then grbp<="111";
	end if;
	if (ll=229 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=243 and ll=229) then grbp<="111";
	end if;
	if (ll=229 and cc>=243 and cc<251) then grbp<="111";
	end if;
	if (cc=49 and ll=230) then grbp<="111";
	end if;
	if (ll=230 and cc>=49 and cc<51) then grbp<="111";
	end if;
	if (ll=230 and cc>=54 and cc<56) then grbp<="111";
	end if;
	if (ll=230 and cc>=104 and cc<112) then grbp<="111";
	end if;
	if (ll=230 and cc>=136 and cc<140) then grbp<="111";
	end if;
	if (ll=230 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (ll=230 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=240 and ll=230) then grbp<="111";
	end if;
	if (cc=243 and ll=230) then grbp<="111";
	end if;
	if (ll=230 and cc>=243 and cc<251) then grbp<="111";
	end if;
	if (cc=54 and ll=231) then grbp<="111";
	end if;
	if (cc=104 and ll=231) then grbp<="111";
	end if;
	if (ll=231 and cc>=104 and cc<112) then grbp<="111";
	end if;
	if (ll=231 and cc>=137 and cc<139) then grbp<="111";
	end if;
	if (ll=231 and cc>=150 and cc<156) then grbp<="111";
	end if;
	if (ll=231 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=239 and ll=231) then grbp<="111";
	end if;
	if (cc=242 and ll=231) then grbp<="111";
	end if;
	if (cc=244 and ll=231) then grbp<="111";
	end if;
	if (ll=231 and cc>=244 and cc<251) then grbp<="111";
	end if;
	if (cc=104 and ll=232) then grbp<="111";
	end if;
	if (ll=232 and cc>=104 and cc<111) then grbp<="111";
	end if;
	if (ll=232 and cc>=150 and cc<156) then grbp<="111";
	end if;
	if (cc=241 and ll=232) then grbp<="111";
	end if;
	if (ll=232 and cc>=241 and cc<243) then grbp<="111";
	end if;
	if (ll=232 and cc>=244 and cc<251) then grbp<="111";
	end if;
	if (ll=233 and cc>=24 and cc<26) then grbp<="111";
	end if;
	if (cc=63 and ll=233) then grbp<="111";
	end if;
	if (cc=103 and ll=233) then grbp<="111";
	end if;
	if (ll=233 and cc>=103 and cc<111) then grbp<="111";
	end if;
	if (ll=233 and cc>=136 and cc<138) then grbp<="111";
	end if;
	if (ll=233 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (ll=233 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (cc=212 and ll=233) then grbp<="111";
	end if;
	if (cc=214 and ll=233) then grbp<="111";
	end if;
	if (cc=240 and ll=233) then grbp<="111";
	end if;
	if (ll=233 and cc>=240 and cc<251) then grbp<="111";
	end if;
	if (ll=234 and cc>=24 and cc<26) then grbp<="111";
	end if;
	if (ll=234 and cc>=47 and cc<49) then grbp<="111";
	end if;
	if (cc=103 and ll=234) then grbp<="111";
	end if;
	if (ll=234 and cc>=103 and cc<110) then grbp<="111";
	end if;
	if (ll=234 and cc>=136 and cc<140) then grbp<="111";
	end if;
	if (ll=234 and cc>=150 and cc<158) then grbp<="111";
	end if;
	if (ll=234 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (cc=216 and ll=234) then grbp<="111";
	end if;
	if (cc=237 and ll=234) then grbp<="111";
	end if;
	if (ll=234 and cc>=237 and cc<251) then grbp<="111";
	end if;
	if (cc=47 and ll=235) then grbp<="111";
	end if;
	if (cc=103 and ll=235) then grbp<="111";
	end if;
	if (ll=235 and cc>=103 and cc<110) then grbp<="111";
	end if;
	if (cc=133 and ll=235) then grbp<="111";
	end if;
	if (ll=235 and cc>=133 and cc<140) then grbp<="111";
	end if;
	if (ll=235 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (ll=235 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (ll=235 and cc>=236 and cc<251) then grbp<="111";
	end if;
	if (ll=236 and cc>=24 and cc<27) then grbp<="111";
	end if;
	if (cc=102 and ll=236) then grbp<="111";
	end if;
	if (ll=236 and cc>=102 and cc<109) then grbp<="111";
	end if;
	if (ll=236 and cc>=121 and cc<126) then grbp<="111";
	end if;
	if (ll=236 and cc>=130 and cc<140) then grbp<="111";
	end if;
	if (ll=236 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (ll=236 and cc>=180 and cc<182) then grbp<="111";
	end if;
	if (ll=236 and cc>=236 and cc<251) then grbp<="111";
	end if;
	if (ll=237 and cc>=23 and cc<26) then grbp<="111";
	end if;
	if (ll=237 and cc>=102 and cc<109) then grbp<="111";
	end if;
	if (ll=237 and cc>=121 and cc<140) then grbp<="111";
	end if;
	if (ll=237 and cc>=150 and cc<158) then grbp<="111";
	end if;
	if (cc=180 and ll=237) then grbp<="111";
	end if;
	if (ll=237 and cc>=180 and cc<183) then grbp<="111";
	end if;
	if (ll=237 and cc>=235 and cc<251) then grbp<="111";
	end if;
	if (cc=24 and ll=238) then grbp<="111";
	end if;
	if (cc=77 and ll=238) then grbp<="111";
	end if;
	if (cc=82 and ll=238) then grbp<="111";
	end if;
	if (cc=102 and ll=238) then grbp<="111";
	end if;
	if (ll=238 and cc>=102 and cc<108) then grbp<="111";
	end if;
	if (ll=238 and cc>=120 and cc<139) then grbp<="111";
	end if;
	if (ll=238 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (ll=238 and cc>=180 and cc<183) then grbp<="111";
	end if;
	if (cc=223 and ll=238) then grbp<="111";
	end if;
	if (cc=235 and ll=238) then grbp<="111";
	end if;
	if (ll=238 and cc>=235 and cc<251) then grbp<="111";
	end if;
	if (cc=25 and ll=239) then grbp<="111";
	end if;
	if (cc=51 and ll=239) then grbp<="111";
	end if;
	if (cc=82 and ll=239) then grbp<="111";
	end if;
	if (cc=101 and ll=239) then grbp<="111";
	end if;
	if (ll=239 and cc>=101 and cc<108) then grbp<="111";
	end if;
	if (ll=239 and cc>=121 and cc<139) then grbp<="111";
	end if;
	if (ll=239 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (ll=239 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (cc=212 and ll=239) then grbp<="111";
	end if;
	if (cc=235 and ll=239) then grbp<="111";
	end if;
	if (ll=239 and cc>=235 and cc<245) then grbp<="111";
	end if;
	if (ll=239 and cc>=247 and cc<251) then grbp<="111";
	end if;
	if (ll=240 and cc>=48 and cc<52) then grbp<="111";
	end if;
	if (cc=101 and ll=240) then grbp<="111";
	end if;
	if (ll=240 and cc>=101 and cc<107) then grbp<="111";
	end if;
	if (ll=240 and cc>=120 and cc<138) then grbp<="111";
	end if;
	if (ll=240 and cc>=150 and cc<159) then grbp<="111";
	end if;
	if (ll=240 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (cc=216 and ll=240) then grbp<="111";
	end if;
	if (cc=234 and ll=240) then grbp<="111";
	end if;
	if (ll=240 and cc>=234 and cc<242) then grbp<="111";
	end if;
	if (ll=240 and cc>=243 and cc<246) then grbp<="111";
	end if;
	if (ll=240 and cc>=247 and cc<251) then grbp<="111";
	end if;
	if (cc=46 and ll=241) then grbp<="111";
	end if;
	if (ll=241 and cc>=46 and cc<49) then grbp<="111";
	end if;
	if (cc=101 and ll=241) then grbp<="111";
	end if;
	if (ll=241 and cc>=101 and cc<107) then grbp<="111";
	end if;
	if (ll=241 and cc>=121 and cc<139) then grbp<="111";
	end if;
	if (ll=241 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=241 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (ll=241 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=241 and cc>=234 and cc<242) then grbp<="111";
	end if;
	if (ll=241 and cc>=243 and cc<251) then grbp<="111";
	end if;
	if (ll=242 and cc>=42 and cc<48) then grbp<="111";
	end if;
	if (ll=242 and cc>=101 and cc<106) then grbp<="111";
	end if;
	if (ll=242 and cc>=121 and cc<138) then grbp<="111";
	end if;
	if (ll=242 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=242 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (cc=233 and ll=242) then grbp<="111";
	end if;
	if (ll=242 and cc>=233 and cc<245) then grbp<="111";
	end if;
	if (ll=242 and cc>=246 and cc<251) then grbp<="111";
	end if;
	if (cc=100 and ll=243) then grbp<="111";
	end if;
	if (ll=243 and cc>=100 and cc<106) then grbp<="111";
	end if;
	if (ll=243 and cc>=121 and cc<139) then grbp<="111";
	end if;
	if (ll=243 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=243 and cc>=181 and cc<184) then grbp<="111";
	end if;
	if (cc=233 and ll=243) then grbp<="111";
	end if;
	if (ll=243 and cc>=233 and cc<242) then grbp<="111";
	end if;
	if (ll=243 and cc>=243 and cc<251) then grbp<="111";
	end if;
	if (cc=100 and ll=244) then grbp<="111";
	end if;
	if (ll=244 and cc>=100 and cc<105) then grbp<="111";
	end if;
	if (ll=244 and cc>=122 and cc<139) then grbp<="111";
	end if;
	if (ll=244 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=244 and cc>=181 and cc<184) then grbp<="111";
	end if;
	if (cc=213 and ll=244) then grbp<="111";
	end if;
	if (cc=233 and ll=244) then grbp<="111";
	end if;
	if (ll=244 and cc>=233 and cc<240) then grbp<="111";
	end if;
	if (cc=245 and ll=244) then grbp<="111";
	end if;
	if (ll=244 and cc>=245 and cc<251) then grbp<="111";
	end if;
	if (cc=100 and ll=245) then grbp<="111";
	end if;
	if (ll=245 and cc>=100 and cc<105) then grbp<="111";
	end if;
	if (ll=245 and cc>=122 and cc<138) then grbp<="111";
	end if;
	if (ll=245 and cc>=151 and cc<161) then grbp<="111";
	end if;
	if (cc=183 and ll=245) then grbp<="111";
	end if;
	if (cc=199 and ll=245) then grbp<="111";
	end if;
	if (cc=210 and ll=245) then grbp<="111";
	end if;
	if (cc=232 and ll=245) then grbp<="111";
	end if;
	if (ll=245 and cc>=232 and cc<237) then grbp<="111";
	end if;
	if (ll=245 and cc>=239 and cc<242) then grbp<="111";
	end if;
	if (ll=245 and cc>=244 and cc<251) then grbp<="111";
	end if;
	if (cc=100 and ll=246) then grbp<="111";
	end if;
	if (ll=246 and cc>=100 and cc<105) then grbp<="111";
	end if;
	if (ll=246 and cc>=123 and cc<138) then grbp<="111";
	end if;
	if (ll=246 and cc>=151 and cc<161) then grbp<="111";
	end if;
	if (cc=183 and ll=246) then grbp<="111";
	end if;
	if (cc=205 and ll=246) then grbp<="111";
	end if;
	if (cc=212 and ll=246) then grbp<="111";
	end if;
	if (cc=231 and ll=246) then grbp<="111";
	end if;
	if (ll=246 and cc>=231 and cc<238) then grbp<="111";
	end if;
	if (ll=246 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (ll=247 and cc>=99 and cc<104) then grbp<="111";
	end if;
	if (ll=247 and cc>=122 and cc<137) then grbp<="111";
	end if;
	if (ll=247 and cc>=151 and cc<161) then grbp<="111";
	end if;
	if (cc=183 and ll=247) then grbp<="111";
	end if;
	if (cc=231 and ll=247) then grbp<="111";
	end if;
	if (ll=247 and cc>=231 and cc<234) then grbp<="111";
	end if;
	if (ll=247 and cc>=235 and cc<238) then grbp<="111";
	end if;
	if (ll=247 and cc>=240 and cc<251) then grbp<="111";
	end if;
	if (ll=248 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (cc=99 and ll=248) then grbp<="111";
	end if;
	if (ll=248 and cc>=99 and cc<104) then grbp<="111";
	end if;
	if (cc=125 and ll=248) then grbp<="111";
	end if;
	if (ll=248 and cc>=125 and cc<137) then grbp<="111";
	end if;
	if (ll=248 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (cc=183 and ll=248) then grbp<="111";
	end if;
	if (cc=205 and ll=248) then grbp<="111";
	end if;
	if (cc=231 and ll=248) then grbp<="111";
	end if;
	if (ll=248 and cc>=231 and cc<238) then grbp<="111";
	end if;
	if (ll=248 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (cc=60 and ll=249) then grbp<="111";
	end if;
	if (cc=99 and ll=249) then grbp<="111";
	end if;
	if (ll=249 and cc>=99 and cc<103) then grbp<="111";
	end if;
	if (ll=249 and cc>=125 and cc<137) then grbp<="111";
	end if;
	if (ll=249 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (cc=199 and ll=249) then grbp<="111";
	end if;
	if (cc=216 and ll=249) then grbp<="111";
	end if;
	if (cc=230 and ll=249) then grbp<="111";
	end if;
	if (cc=232 and ll=249) then grbp<="111";
	end if;
	if (ll=249 and cc>=232 and cc<236) then grbp<="111";
	end if;
	if (ll=249 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (ll=250 and cc>=98 and cc<103) then grbp<="111";
	end if;
	if (ll=250 and cc>=125 and cc<136) then grbp<="111";
	end if;
	if (ll=250 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=250 and cc>=181 and cc<184) then grbp<="111";
	end if;
	if (ll=250 and cc>=197 and cc<199) then grbp<="111";
	end if;
	if (ll=250 and cc>=230 and cc<236) then grbp<="111";
	end if;
	if (cc=240 and ll=250) then grbp<="111";
	end if;
	if (ll=250 and cc>=240 and cc<251) then grbp<="111";
	end if;
	if (cc=86 and ll=251) then grbp<="111";
	end if;
	if (cc=98 and ll=251) then grbp<="111";
	end if;
	if (ll=251 and cc>=98 and cc<103) then grbp<="111";
	end if;
	if (ll=251 and cc>=124 and cc<136) then grbp<="111";
	end if;
	if (ll=251 and cc>=151 and cc<160) then grbp<="111";
	end if;
	if (ll=251 and cc>=181 and cc<184) then grbp<="111";
	end if;
	if (ll=251 and cc>=198 and cc<200) then grbp<="111";
	end if;
	if (ll=251 and cc>=230 and cc<236) then grbp<="111";
	end if;
	if (cc=239 and ll=251) then grbp<="111";
	end if;
	if (ll=251 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (cc=98 and ll=252) then grbp<="111";
	end if;
	if (ll=252 and cc>=98 and cc<102) then grbp<="111";
	end if;
	if (ll=252 and cc>=125 and cc<136) then grbp<="111";
	end if;
	if (ll=252 and cc>=152 and cc<160) then grbp<="111";
	end if;
	if (ll=252 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (cc=233 and ll=252) then grbp<="111";
	end if;
	if (ll=252 and cc>=233 and cc<235) then grbp<="111";
	end if;
	if (ll=252 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (cc=88 and ll=253) then grbp<="111";
	end if;
	if (cc=98 and ll=253) then grbp<="111";
	end if;
	if (ll=253 and cc>=98 and cc<102) then grbp<="111";
	end if;
	if (ll=253 and cc>=125 and cc<136) then grbp<="111";
	end if;
	if (ll=253 and cc>=151 and cc<158) then grbp<="111";
	end if;
	if (cc=181 and ll=253) then grbp<="111";
	end if;
	if (ll=253 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (ll=253 and cc>=230 and cc<233) then grbp<="111";
	end if;
	if (cc=239 and ll=253) then grbp<="111";
	end if;
	if (ll=253 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (cc=41 and ll=254) then grbp<="111";
	end if;
	if (ll=254 and cc>=41 and cc<43) then grbp<="111";
	end if;
	if (cc=63 and ll=254) then grbp<="111";
	end if;
	if (cc=83 and ll=254) then grbp<="111";
	end if;
	if (cc=97 and ll=254) then grbp<="111";
	end if;
	if (ll=254 and cc>=97 and cc<101) then grbp<="111";
	end if;
	if (ll=254 and cc>=123 and cc<125) then grbp<="111";
	end if;
	if (ll=254 and cc>=126 and cc<135) then grbp<="111";
	end if;
	if (cc=151 and ll=254) then grbp<="111";
	end if;
	if (ll=254 and cc>=151 and cc<159) then grbp<="111";
	end if;
	if (ll=254 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (ll=254 and cc>=230 and cc<232) then grbp<="111";
	end if;
	if (ll=254 and cc>=239 and cc<251) then grbp<="111";
	end if;
	if (cc=40 and ll=255) then grbp<="111";
	end if;
	if (cc=83 and ll=255) then grbp<="111";
	end if;
	if (ll=255 and cc>=83 and cc<85) then grbp<="111";
	end if;
	if (ll=255 and cc>=97 and cc<101) then grbp<="111";
	end if;
	if (ll=255 and cc>=125 and cc<137) then grbp<="111";
	end if;
	if (ll=255 and cc>=151 and cc<159) then grbp<="111";
	end if;
	if (ll=255 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (ll=255 and cc>=230 and cc<232) then grbp<="111";
	end if;
	if (cc=237 and ll=255) then grbp<="111";
	end if;
	if (ll=255 and cc>=237 and cc<251) then grbp<="111";
	end if;
	if (cc=83 and ll=256) then grbp<="111";
	end if;
	if (ll=256 and cc>=83 and cc<85) then grbp<="111";
	end if;
	if (ll=256 and cc>=97 and cc<101) then grbp<="111";
	end if;
	if (ll=256 and cc>=128 and cc<135) then grbp<="111";
	end if;
	if (ll=256 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=181 and ll=256) then grbp<="111";
	end if;
	if (ll=256 and cc>=181 and cc<183) then grbp<="111";
	end if;
	if (ll=256 and cc>=229 and cc<232) then grbp<="111";
	end if;
	if (cc=237 and ll=256) then grbp<="111";
	end if;
	if (ll=256 and cc>=237 and cc<251) then grbp<="111";
	end if;
	if (cc=83 and ll=257) then grbp<="111";
	end if;
	if (ll=257 and cc>=83 and cc<86) then grbp<="111";
	end if;
	if (ll=257 and cc>=97 and cc<100) then grbp<="111";
	end if;
	if (cc=132 and ll=257) then grbp<="111";
	end if;
	if (ll=257 and cc>=132 and cc<135) then grbp<="111";
	end if;
	if (ll=257 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=182 and ll=257) then grbp<="111";
	end if;
	if (cc=229 and ll=257) then grbp<="111";
	end if;
	if (ll=257 and cc>=229 and cc<232) then grbp<="111";
	end if;
	if (ll=257 and cc>=234 and cc<251) then grbp<="111";
	end if;
	if (cc=21 and ll=258) then grbp<="111";
	end if;
	if (cc=62 and ll=258) then grbp<="111";
	end if;
	if (cc=84 and ll=258) then grbp<="111";
	end if;
	if (ll=258 and cc>=84 and cc<86) then grbp<="111";
	end if;
	if (ll=258 and cc>=96 and cc<100) then grbp<="111";
	end if;
	if (cc=132 and ll=258) then grbp<="111";
	end if;
	if (ll=258 and cc>=132 and cc<134) then grbp<="111";
	end if;
	if (ll=258 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=182 and ll=258) then grbp<="111";
	end if;
	if (cc=184 and ll=258) then grbp<="111";
	end if;
	if (cc=214 and ll=258) then grbp<="111";
	end if;
	if (cc=229 and ll=258) then grbp<="111";
	end if;
	if (ll=258 and cc>=229 and cc<232) then grbp<="111";
	end if;
	if (ll=258 and cc>=235 and cc<251) then grbp<="111";
	end if;
	if (cc=96 and ll=259) then grbp<="111";
	end if;
	if (ll=259 and cc>=96 and cc<99) then grbp<="111";
	end if;
	if (ll=259 and cc>=129 and cc<132) then grbp<="111";
	end if;
	if (ll=259 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=182 and ll=259) then grbp<="111";
	end if;
	if (cc=227 and ll=259) then grbp<="111";
	end if;
	if (cc=229 and ll=259) then grbp<="111";
	end if;
	if (cc=234 and ll=259) then grbp<="111";
	end if;
	if (cc=236 and ll=259) then grbp<="111";
	end if;
	if (ll=259 and cc>=236 and cc<251) then grbp<="111";
	end if;
	if (cc=96 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=96 and cc<99) then grbp<="111";
	end if;
	if (cc=133 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=133 and cc<135) then grbp<="111";
	end if;
	if (ll=260 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=184 and ll=260) then grbp<="111";
	end if;
	if (cc=196 and ll=260) then grbp<="111";
	end if;
	if (cc=209 and ll=260) then grbp<="111";
	end if;
	if (cc=227 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=227 and cc<231) then grbp<="111";
	end if;
	if (cc=234 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=234 and cc<251) then grbp<="111";
	end if;
	if (cc=96 and ll=261) then grbp<="111";
	end if;
	if (ll=261 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=261 and cc>=130 and cc<135) then grbp<="111";
	end if;
	if (ll=261 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (cc=184 and ll=261) then grbp<="111";
	end if;
	if (cc=227 and ll=261) then grbp<="111";
	end if;
	if (ll=261 and cc>=227 and cc<231) then grbp<="111";
	end if;
	if (ll=261 and cc>=233 and cc<251) then grbp<="111";
	end if;
	if (cc=96 and ll=262) then grbp<="111";
	end if;
	if (cc=130 and ll=262) then grbp<="111";
	end if;
	if (cc=133 and ll=262) then grbp<="111";
	end if;
	if (cc=152 and ll=262) then grbp<="111";
	end if;
	if (ll=262 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (ll=262 and cc>=182 and cc<185) then grbp<="111";
	end if;
	if (cc=227 and ll=262) then grbp<="111";
	end if;
	if (ll=262 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=234 and ll=262) then grbp<="111";
	end if;
	if (ll=262 and cc>=234 and cc<251) then grbp<="111";
	end if;
	if (cc=62 and ll=263) then grbp<="111";
	end if;
	if (cc=91 and ll=263) then grbp<="111";
	end if;
	if (cc=97 and ll=263) then grbp<="111";
	end if;
	if (cc=132 and ll=263) then grbp<="111";
	end if;
	if (cc=152 and ll=263) then grbp<="111";
	end if;
	if (ll=263 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (ll=263 and cc>=182 and cc<184) then grbp<="111";
	end if;
	if (cc=227 and ll=263) then grbp<="111";
	end if;
	if (ll=263 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=263 and cc>=234 and cc<251) then grbp<="111";
	end if;
	if (cc=62 and ll=264) then grbp<="111";
	end if;
	if (cc=90 and ll=264) then grbp<="111";
	end if;
	if (ll=264 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (cc=96 and ll=264) then grbp<="111";
	end if;
	if (ll=264 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=264 and cc>=152 and cc<157) then grbp<="111";
	end if;
	if (ll=264 and cc>=182 and cc<184) then grbp<="111";
	end if;
	if (ll=264 and cc>=197 and cc<199) then grbp<="111";
	end if;
	if (cc=212 and ll=264) then grbp<="111";
	end if;
	if (cc=227 and ll=264) then grbp<="111";
	end if;
	if (ll=264 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (cc=234 and ll=264) then grbp<="111";
	end if;
	if (ll=264 and cc>=234 and cc<251) then grbp<="111";
	end if;
	if (cc=65 and ll=265) then grbp<="111";
	end if;
	if (cc=90 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=90 and cc<97) then grbp<="111";
	end if;
	if (cc=153 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=153 and cc<157) then grbp<="111";
	end if;
	if (ll=265 and cc>=182 and cc<184) then grbp<="111";
	end if;
	if (cc=226 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=233 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=233 and cc<251) then grbp<="111";
	end if;
	if (cc=90 and ll=266) then grbp<="111";
	end if;
	if (ll=266 and cc>=90 and cc<97) then grbp<="111";
	end if;
	if (ll=266 and cc>=153 and cc<157) then grbp<="111";
	end if;
	if (ll=266 and cc>=182 and cc<184) then grbp<="111";
	end if;
	if (cc=225 and ll=266) then grbp<="111";
	end if;
	if (ll=266 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=232 and ll=266) then grbp<="111";
	end if;
	if (ll=266 and cc>=232 and cc<251) then grbp<="111";
	end if;
	if (cc=54 and ll=267) then grbp<="111";
	end if;
	if (cc=62 and ll=267) then grbp<="111";
	end if;
	if (ll=267 and cc>=62 and cc<64) then grbp<="111";
	end if;
	if (ll=267 and cc>=89 and cc<96) then grbp<="111";
	end if;
	if (cc=153 and ll=267) then grbp<="111";
	end if;
	if (ll=267 and cc>=153 and cc<157) then grbp<="111";
	end if;
	if (ll=267 and cc>=182 and cc<184) then grbp<="111";
	end if;
	if (cc=226 and ll=267) then grbp<="111";
	end if;
	if (ll=267 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=232 and ll=267) then grbp<="111";
	end if;
	if (ll=267 and cc>=232 and cc<251) then grbp<="111";
	end if;
	if (ll=268 and cc>=20 and cc<23) then grbp<="111";
	end if;
	if (cc=62 and ll=268) then grbp<="111";
	end if;
	if (ll=268 and cc>=62 and cc<64) then grbp<="111";
	end if;
	if (cc=89 and ll=268) then grbp<="111";
	end if;
	if (ll=268 and cc>=89 and cc<96) then grbp<="111";
	end if;
	if (ll=268 and cc>=153 and cc<157) then grbp<="111";
	end if;
	if (cc=195 and ll=268) then grbp<="111";
	end if;
	if (cc=225 and ll=268) then grbp<="111";
	end if;
	if (cc=228 and ll=268) then grbp<="111";
	end if;
	if (cc=232 and ll=268) then grbp<="111";
	end if;
	if (ll=268 and cc>=232 and cc<251) then grbp<="111";
	end if;
	if (cc=63 and ll=269) then grbp<="111";
	end if;
	if (cc=80 and ll=269) then grbp<="111";
	end if;
	if (cc=89 and ll=269) then grbp<="111";
	end if;
	if (ll=269 and cc>=89 and cc<96) then grbp<="111";
	end if;
	if (ll=269 and cc>=154 and cc<158) then grbp<="111";
	end if;
	if (cc=185 and ll=269) then grbp<="111";
	end if;
	if (cc=227 and ll=269) then grbp<="111";
	end if;
	if (ll=269 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=269 and cc>=230 and cc<251) then grbp<="111";
	end if;
	if (cc=63 and ll=270) then grbp<="111";
	end if;
	if (cc=90 and ll=270) then grbp<="111";
	end if;
	if (ll=270 and cc>=90 and cc<95) then grbp<="111";
	end if;
	if (ll=270 and cc>=154 and cc<157) then grbp<="111";
	end if;
	if (cc=185 and ll=270) then grbp<="111";
	end if;
	if (cc=226 and ll=270) then grbp<="111";
	end if;
	if (ll=270 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=270 and cc>=229 and cc<251) then grbp<="111";
	end if;
	if (ll=271 and cc>=20 and cc<22) then grbp<="111";
	end if;
	if (cc=66 and ll=271) then grbp<="111";
	end if;
	if (cc=92 and ll=271) then grbp<="111";
	end if;
	if (ll=271 and cc>=92 and cc<94) then grbp<="111";
	end if;
	if (ll=271 and cc>=153 and cc<157) then grbp<="111";
	end if;
	if (cc=226 and ll=271) then grbp<="111";
	end if;
	if (ll=271 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=271 and cc>=230 and cc<251) then grbp<="111";
	end if;
	if (cc=66 and ll=272) then grbp<="111";
	end if;
	if (cc=92 and ll=272) then grbp<="111";
	end if;
	if (ll=272 and cc>=92 and cc<94) then grbp<="111";
	end if;
	if (cc=152 and ll=272) then grbp<="111";
	end if;
	if (ll=272 and cc>=152 and cc<158) then grbp<="111";
	end if;
	if (cc=226 and ll=272) then grbp<="111";
	end if;
	if (cc=230 and ll=272) then grbp<="111";
	end if;
	if (ll=272 and cc>=230 and cc<251) then grbp<="111";
	end if;
	if (ll=273 and cc>=24 and cc<27) then grbp<="111";
	end if;
	if (cc=87 and ll=273) then grbp<="111";
	end if;
	if (cc=92 and ll=273) then grbp<="111";
	end if;
	if (ll=273 and cc>=92 and cc<94) then grbp<="111";
	end if;
	if (cc=151 and ll=273) then grbp<="111";
	end if;
	if (ll=273 and cc>=151 and cc<157) then grbp<="111";
	end if;
	if (cc=207 and ll=273) then grbp<="111";
	end if;
	if (cc=225 and ll=273) then grbp<="111";
	end if;
	if (cc=227 and ll=273) then grbp<="111";
	end if;
	if (cc=229 and ll=273) then grbp<="111";
	end if;
	if (ll=273 and cc>=229 and cc<251) then grbp<="111";
	end if;
	if (cc=86 and ll=274) then grbp<="111";
	end if;
	if (ll=274 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (cc=135 and ll=274) then grbp<="111";
	end if;
	if (cc=150 and ll=274) then grbp<="111";
	end if;
	if (ll=274 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (cc=226 and ll=274) then grbp<="111";
	end if;
	if (cc=228 and ll=274) then grbp<="111";
	end if;
	if (ll=274 and cc>=228 and cc<251) then grbp<="111";
	end if;
	if (cc=66 and ll=275) then grbp<="111";
	end if;
	if (cc=85 and ll=275) then grbp<="111";
	end if;
	if (ll=275 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=275 and cc>=91 and cc<93) then grbp<="111";
	end if;
	if (cc=150 and ll=275) then grbp<="111";
	end if;
	if (ll=275 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (ll=275 and cc>=183 and cc<185) then grbp<="111";
	end if;
	if (cc=228 and ll=275) then grbp<="111";
	end if;
	if (ll=275 and cc>=228 and cc<251) then grbp<="111";
	end if;
	if (cc=66 and ll=276) then grbp<="111";
	end if;
	if (cc=84 and ll=276) then grbp<="111";
	end if;
	if (ll=276 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=276 and cc>=91 and cc<93) then grbp<="111";
	end if;
	if (ll=276 and cc>=147 and cc<149) then grbp<="111";
	end if;
	if (ll=276 and cc>=150 and cc<157) then grbp<="111";
	end if;
	if (ll=276 and cc>=183 and cc<185) then grbp<="111";
	end if;
	if (ll=276 and cc>=229 and cc<251) then grbp<="111";
	end if;
	if (ll=277 and cc>=23 and cc<25) then grbp<="111";
	end if;
	if (cc=83 and ll=277) then grbp<="111";
	end if;
	if (ll=277 and cc>=83 and cc<86) then grbp<="111";
	end if;
	if (ll=277 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (ll=277 and cc>=146 and cc<156) then grbp<="111";
	end if;
	if (ll=277 and cc>=183 and cc<185) then grbp<="111";
	end if;
	if (cc=228 and ll=277) then grbp<="111";
	end if;
	if (ll=277 and cc>=228 and cc<251) then grbp<="111";
	end if;
	if (cc=83 and ll=278) then grbp<="111";
	end if;
	if (ll=278 and cc>=83 and cc<86) then grbp<="111";
	end if;
	if (ll=278 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (cc=146 and ll=278) then grbp<="111";
	end if;
	if (ll=278 and cc>=146 and cc<157) then grbp<="111";
	end if;
	if (ll=278 and cc>=183 and cc<185) then grbp<="111";
	end if;
	if (cc=228 and ll=278) then grbp<="111";
	end if;
	if (ll=278 and cc>=228 and cc<251) then grbp<="111";
	end if;
	if (cc=82 and ll=279) then grbp<="111";
	end if;
	if (ll=279 and cc>=82 and cc<86) then grbp<="111";
	end if;
	if (cc=146 and ll=279) then grbp<="111";
	end if;
	if (ll=279 and cc>=146 and cc<157) then grbp<="111";
	end if;
	if (cc=228 and ll=279) then grbp<="111";
	end if;
	if (ll=279 and cc>=228 and cc<251) then grbp<="111";
	end if;
	if (ll=280 and cc>=24 and cc<26) then grbp<="111";
	end if;
	if (cc=80 and ll=280) then grbp<="111";
	end if;
	if (cc=82 and ll=280) then grbp<="111";
	end if;
	if (ll=280 and cc>=82 and cc<85) then grbp<="111";
	end if;
	if (cc=145 and ll=280) then grbp<="111";
	end if;
	if (ll=280 and cc>=145 and cc<156) then grbp<="111";
	end if;
	if (cc=227 and ll=280) then grbp<="111";
	end if;
	if (ll=280 and cc>=227 and cc<251) then grbp<="111";
	end if;
	if (cc=81 and ll=281) then grbp<="111";
	end if;
	if (ll=281 and cc>=81 and cc<85) then grbp<="111";
	end if;
	if (cc=145 and ll=281) then grbp<="111";
	end if;
	if (ll=281 and cc>=145 and cc<157) then grbp<="111";
	end if;
	if (cc=227 and ll=281) then grbp<="111";
	end if;
	if (ll=281 and cc>=227 and cc<251) then grbp<="111";
	end if;
	if (cc=81 and ll=282) then grbp<="111";
	end if;
	if (ll=282 and cc>=81 and cc<85) then grbp<="111";
	end if;
	if (cc=145 and ll=282) then grbp<="111";
	end if;
	if (ll=282 and cc>=145 and cc<156) then grbp<="111";
	end if;
	if (cc=224 and ll=282) then grbp<="111";
	end if;
	if (ll=282 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (ll=282 and cc>=227 and cc<251) then grbp<="111";
	end if;
	if (ll=283 and cc>=81 and cc<84) then grbp<="111";
	end if;
	if (cc=144 and ll=283) then grbp<="111";
	end if;
	if (ll=283 and cc>=144 and cc<156) then grbp<="111";
	end if;
	if (cc=227 and ll=283) then grbp<="111";
	end if;
	if (ll=283 and cc>=227 and cc<251) then grbp<="111";
	end if;
	if (ll=284 and cc>=24 and cc<26) then grbp<="111";
	end if;
	if (cc=81 and ll=284) then grbp<="111";
	end if;
	if (ll=284 and cc>=81 and cc<84) then grbp<="111";
	end if;
	if (cc=145 and ll=284) then grbp<="111";
	end if;
	if (ll=284 and cc>=145 and cc<156) then grbp<="111";
	end if;
	if (cc=206 and ll=284) then grbp<="111";
	end if;
	if (cc=226 and ll=284) then grbp<="111";
	end if;
	if (ll=284 and cc>=226 and cc<251) then grbp<="111";
	end if;
	if (ll=285 and cc>=24 and cc<26) then grbp<="111";
	end if;
	if (cc=69 and ll=285) then grbp<="111";
	end if;
	if (cc=80 and ll=285) then grbp<="111";
	end if;
	if (ll=285 and cc>=80 and cc<83) then grbp<="111";
	end if;
	if (cc=144 and ll=285) then grbp<="111";
	end if;
	if (ll=285 and cc>=144 and cc<156) then grbp<="111";
	end if;
	if (cc=225 and ll=285) then grbp<="111";
	end if;
	if (ll=285 and cc>=225 and cc<251) then grbp<="111";
	end if;
	if (cc=69 and ll=286) then grbp<="111";
	end if;
	if (cc=76 and ll=286) then grbp<="111";
	end if;
	if (ll=286 and cc>=76 and cc<83) then grbp<="111";
	end if;
	if (cc=148 and ll=286) then grbp<="111";
	end if;
	if (ll=286 and cc>=148 and cc<156) then grbp<="111";
	end if;
	if (cc=226 and ll=286) then grbp<="111";
	end if;
	if (ll=286 and cc>=226 and cc<251) then grbp<="111";
	end if;
	if (cc=77 and ll=287) then grbp<="111";
	end if;
	if (ll=287 and cc>=77 and cc<82) then grbp<="111";
	end if;
	if (cc=150 and ll=287) then grbp<="111";
	end if;
	if (cc=184 and ll=287) then grbp<="111";
	end if;
	if (cc=225 and ll=287) then grbp<="111";
	end if;
	if (ll=287 and cc>=225 and cc<251) then grbp<="111";
	end if;
	if (cc=26 and ll=288) then grbp<="111";
	end if;
	if (cc=76 and ll=288) then grbp<="111";
	end if;
	if (ll=288 and cc>=76 and cc<82) then grbp<="111";
	end if;
	if (cc=184 and ll=288) then grbp<="111";
	end if;
	if (cc=224 and ll=288) then grbp<="111";
	end if;
	if (ll=288 and cc>=224 and cc<251) then grbp<="111";
	end if;
	if (cc=21 and ll=289) then grbp<="111";
	end if;
	if (ll=289 and cc>=21 and cc<23) then grbp<="111";
	end if;
	if (cc=76 and ll=289) then grbp<="111";
	end if;
	if (ll=289 and cc>=76 and cc<81) then grbp<="111";
	end if;
	if (cc=184 and ll=289) then grbp<="111";
	end if;
	if (cc=224 and ll=289) then grbp<="111";
	end if;
	if (ll=289 and cc>=224 and cc<251) then grbp<="111";
	end if;
	if (cc=41 and ll=290) then grbp<="111";
	end if;
	if (cc=73 and ll=290) then grbp<="111";
	end if;
	if (ll=290 and cc>=73 and cc<75) then grbp<="111";
	end if;
	if (ll=290 and cc>=76 and cc<81) then grbp<="111";
	end if;
	if (cc=184 and ll=290) then grbp<="111";
	end if;
	if (cc=225 and ll=290) then grbp<="111";
	end if;
	if (ll=290 and cc>=225 and cc<251) then grbp<="111";
	end if;
	if (cc=76 and ll=291) then grbp<="111";
	end if;
	if (ll=291 and cc>=76 and cc<81) then grbp<="111";
	end if;
	if (cc=184 and ll=291) then grbp<="111";
	end if;
	if (cc=194 and ll=291) then grbp<="111";
	end if;
	if (cc=224 and ll=291) then grbp<="111";
	end if;
	if (ll=291 and cc>=224 and cc<251) then grbp<="111";
	end if;
	if (cc=21 and ll=292) then grbp<="111";
	end if;
	if (cc=67 and ll=292) then grbp<="111";
	end if;
	if (cc=76 and ll=292) then grbp<="111";
	end if;
	if (ll=292 and cc>=76 and cc<80) then grbp<="111";
	end if;
	if (cc=184 and ll=292) then grbp<="111";
	end if;
	if (cc=223 and ll=292) then grbp<="111";
	end if;
	if (ll=292 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=24 and ll=293) then grbp<="111";
	end if;
	if (cc=26 and ll=293) then grbp<="111";
	end if;
	if (cc=77 and ll=293) then grbp<="111";
	end if;
	if (ll=293 and cc>=77 and cc<80) then grbp<="111";
	end if;
	if (cc=205 and ll=293) then grbp<="111";
	end if;
	if (cc=209 and ll=293) then grbp<="111";
	end if;
	if (cc=211 and ll=293) then grbp<="111";
	end if;
	if (cc=223 and ll=293) then grbp<="111";
	end if;
	if (ll=293 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=24 and ll=294) then grbp<="111";
	end if;
	if (cc=26 and ll=294) then grbp<="111";
	end if;
	if (cc=33 and ll=294) then grbp<="111";
	end if;
	if (cc=57 and ll=294) then grbp<="111";
	end if;
	if (cc=77 and ll=294) then grbp<="111";
	end if;
	if (ll=294 and cc>=77 and cc<80) then grbp<="111";
	end if;
	if (cc=147 and ll=294) then grbp<="111";
	end if;
	if (ll=294 and cc>=147 and cc<151) then grbp<="111";
	end if;
	if (cc=223 and ll=294) then grbp<="111";
	end if;
	if (ll=294 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=57 and ll=295) then grbp<="111";
	end if;
	if (cc=77 and ll=295) then grbp<="111";
	end if;
	if (ll=295 and cc>=77 and cc<79) then grbp<="111";
	end if;
	if (ll=295 and cc>=83 and cc<85) then grbp<="111";
	end if;
	if (ll=295 and cc>=143 and cc<151) then grbp<="111";
	end if;
	if (cc=223 and ll=295) then grbp<="111";
	end if;
	if (ll=295 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=23 and ll=296) then grbp<="111";
	end if;
	if (cc=57 and ll=296) then grbp<="111";
	end if;
	if (cc=77 and ll=296) then grbp<="111";
	end if;
	if (ll=296 and cc>=77 and cc<79) then grbp<="111";
	end if;
	if (cc=143 and ll=296) then grbp<="111";
	end if;
	if (ll=296 and cc>=143 and cc<151) then grbp<="111";
	end if;
	if (ll=296 and cc>=184 and cc<186) then grbp<="111";
	end if;
	if (ll=296 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=29 and ll=297) then grbp<="111";
	end if;
	if (cc=57 and ll=297) then grbp<="111";
	end if;
	if (cc=77 and ll=297) then grbp<="111";
	end if;
	if (cc=83 and ll=297) then grbp<="111";
	end if;
	if (cc=145 and ll=297) then grbp<="111";
	end if;
	if (cc=149 and ll=297) then grbp<="111";
	end if;
	if (ll=297 and cc>=149 and cc<151) then grbp<="111";
	end if;
	if (cc=223 and ll=297) then grbp<="111";
	end if;
	if (ll=297 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=27 and ll=298) then grbp<="111";
	end if;
	if (ll=298 and cc>=27 and cc<31) then grbp<="111";
	end if;
	if (cc=45 and ll=298) then grbp<="111";
	end if;
	if (cc=56 and ll=298) then grbp<="111";
	end if;
	if (ll=298 and cc>=56 and cc<58) then grbp<="111";
	end if;
	if (ll=298 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=298) then grbp<="111";
	end if;
	if (cc=223 and ll=298) then grbp<="111";
	end if;
	if (ll=298 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (ll=299 and cc>=25 and cc<31) then grbp<="111";
	end if;
	if (cc=71 and ll=299) then grbp<="111";
	end if;
	if (cc=76 and ll=299) then grbp<="111";
	end if;
	if (ll=299 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (ll=299 and cc>=81 and cc<83) then grbp<="111";
	end if;
	if (cc=187 and ll=299) then grbp<="111";
	end if;
	if (cc=223 and ll=299) then grbp<="111";
	end if;
	if (ll=299 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (ll=300 and cc>=26 and cc<29) then grbp<="111";
	end if;
	if (cc=56 and ll=300) then grbp<="111";
	end if;
	if (cc=71 and ll=300) then grbp<="111";
	end if;
	if (ll=300 and cc>=71 and cc<73) then grbp<="111";
	end if;
	if (ll=300 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=300) then grbp<="111";
	end if;
	if (cc=187 and ll=300) then grbp<="111";
	end if;
	if (cc=223 and ll=300) then grbp<="111";
	end if;
	if (ll=300 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=22 and ll=301) then grbp<="111";
	end if;
	if (cc=26 and ll=301) then grbp<="111";
	end if;
	if (cc=56 and ll=301) then grbp<="111";
	end if;
	if (cc=59 and ll=301) then grbp<="111";
	end if;
	if (cc=72 and ll=301) then grbp<="111";
	end if;
	if (cc=76 and ll=301) then grbp<="111";
	end if;
	if (ll=301 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=301) then grbp<="111";
	end if;
	if (cc=187 and ll=301) then grbp<="111";
	end if;
	if (cc=222 and ll=301) then grbp<="111";
	end if;
	if (ll=301 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=26 and ll=302) then grbp<="111";
	end if;
	if (cc=36 and ll=302) then grbp<="111";
	end if;
	if (cc=56 and ll=302) then grbp<="111";
	end if;
	if (cc=72 and ll=302) then grbp<="111";
	end if;
	if (cc=76 and ll=302) then grbp<="111";
	end if;
	if (ll=302 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=302) then grbp<="111";
	end if;
	if (cc=187 and ll=302) then grbp<="111";
	end if;
	if (cc=223 and ll=302) then grbp<="111";
	end if;
	if (ll=302 and cc>=223 and cc<251) then grbp<="111";
	end if;
	if (cc=36 and ll=303) then grbp<="111";
	end if;
	if (cc=56 and ll=303) then grbp<="111";
	end if;
	if (cc=67 and ll=303) then grbp<="111";
	end if;
	if (cc=76 and ll=303) then grbp<="111";
	end if;
	if (ll=303 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=303) then grbp<="111";
	end if;
	if (cc=187 and ll=303) then grbp<="111";
	end if;
	if (cc=222 and ll=303) then grbp<="111";
	end if;
	if (ll=303 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=36 and ll=304) then grbp<="111";
	end if;
	if (cc=56 and ll=304) then grbp<="111";
	end if;
	if (ll=304 and cc>=56 and cc<58) then grbp<="111";
	end if;
	if (cc=76 and ll=304) then grbp<="111";
	end if;
	if (cc=79 and ll=304) then grbp<="111";
	end if;
	if (cc=185 and ll=304) then grbp<="111";
	end if;
	if (cc=187 and ll=304) then grbp<="111";
	end if;
	if (cc=207 and ll=304) then grbp<="111";
	end if;
	if (cc=222 and ll=304) then grbp<="111";
	end if;
	if (ll=304 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=55 and ll=305) then grbp<="111";
	end if;
	if (ll=305 and cc>=55 and cc<58) then grbp<="111";
	end if;
	if (cc=76 and ll=305) then grbp<="111";
	end if;
	if (ll=305 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=185 and ll=305) then grbp<="111";
	end if;
	if (cc=187 and ll=305) then grbp<="111";
	end if;
	if (cc=222 and ll=305) then grbp<="111";
	end if;
	if (ll=305 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=55 and ll=306) then grbp<="111";
	end if;
	if (ll=306 and cc>=55 and cc<57) then grbp<="111";
	end if;
	if (ll=306 and cc>=76 and cc<79) then grbp<="111";
	end if;
	if (ll=306 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=222 and ll=306) then grbp<="111";
	end if;
	if (ll=306 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=25 and ll=307) then grbp<="111";
	end if;
	if (ll=307 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (ll=307 and cc>=55 and cc<57) then grbp<="111";
	end if;
	if (cc=75 and ll=307) then grbp<="111";
	end if;
	if (ll=307 and cc>=75 and cc<79) then grbp<="111";
	end if;
	if (ll=307 and cc>=142 and cc<144) then grbp<="111";
	end if;
	if (cc=185 and ll=307) then grbp<="111";
	end if;
	if (ll=307 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=222 and ll=307) then grbp<="111";
	end if;
	if (ll=307 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=61 and ll=308) then grbp<="111";
	end if;
	if (cc=75 and ll=308) then grbp<="111";
	end if;
	if (ll=308 and cc>=75 and cc<78) then grbp<="111";
	end if;
	if (ll=308 and cc>=141 and cc<145) then grbp<="111";
	end if;
	if (ll=308 and cc>=185 and cc<188) then grbp<="111";
	end if;
	if (cc=198 and ll=308) then grbp<="111";
	end if;
	if (cc=204 and ll=308) then grbp<="111";
	end if;
	if (cc=209 and ll=308) then grbp<="111";
	end if;
	if (cc=222 and ll=308) then grbp<="111";
	end if;
	if (ll=308 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=76 and ll=309) then grbp<="111";
	end if;
	if (ll=309 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (ll=309 and cc>=141 and cc<146) then grbp<="111";
	end if;
	if (cc=185 and ll=309) then grbp<="111";
	end if;
	if (ll=309 and cc>=185 and cc<188) then grbp<="111";
	end if;
	if (cc=199 and ll=309) then grbp<="111";
	end if;
	if (cc=204 and ll=309) then grbp<="111";
	end if;
	if (cc=222 and ll=309) then grbp<="111";
	end if;
	if (ll=309 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (ll=310 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (ll=310 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (ll=310 and cc>=140 and cc<149) then grbp<="111";
	end if;
	if (ll=310 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=197 and ll=310) then grbp<="111";
	end if;
	if (cc=222 and ll=310) then grbp<="111";
	end if;
	if (ll=310 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=137 and ll=311) then grbp<="111";
	end if;
	if (ll=311 and cc>=137 and cc<139) then grbp<="111";
	end if;
	if (ll=311 and cc>=140 and cc<149) then grbp<="111";
	end if;
	if (ll=311 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (ll=311 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (cc=26 and ll=312) then grbp<="111";
	end if;
	if (cc=69 and ll=312) then grbp<="111";
	end if;
	if (cc=76 and ll=312) then grbp<="111";
	end if;
	if (cc=136 and ll=312) then grbp<="111";
	end if;
	if (ll=312 and cc>=136 and cc<149) then grbp<="111";
	end if;
	if (ll=312 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=195 and ll=312) then grbp<="111";
	end if;
	if (cc=200 and ll=312) then grbp<="111";
	end if;
	if (cc=209 and ll=312) then grbp<="111";
	end if;
	if (cc=221 and ll=312) then grbp<="111";
	end if;
	if (ll=312 and cc>=221 and cc<251) then grbp<="111";
	end if;
	if (cc=63 and ll=313) then grbp<="111";
	end if;
	if (cc=69 and ll=313) then grbp<="111";
	end if;
	if (cc=137 and ll=313) then grbp<="111";
	end if;
	if (ll=313 and cc>=137 and cc<149) then grbp<="111";
	end if;
	if (ll=313 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=200 and ll=313) then grbp<="111";
	end if;
	if (cc=222 and ll=313) then grbp<="111";
	end if;
	if (ll=313 and cc>=222 and cc<251) then grbp<="111";
	end if;
	if (ll=314 and cc>=137 and cc<149) then grbp<="111";
	end if;
	if (ll=314 and cc>=185 and cc<187) then grbp<="111";
	end if;
	if (cc=199 and ll=314) then grbp<="111";
	end if;
	if (cc=221 and ll=314) then grbp<="111";
	end if;
	if (ll=314 and cc>=221 and cc<251) then grbp<="111";
	end if;
	if (ll=315 and cc>=138 and cc<149) then grbp<="111";
	end if;
	if (cc=200 and ll=315) then grbp<="111";
	end if;
	if (cc=221 and ll=315) then grbp<="111";
	end if;
	if (ll=315 and cc>=221 and cc<249) then grbp<="111";
	end if;
	if (cc=66 and ll=316) then grbp<="111";
	end if;
	if (cc=138 and ll=316) then grbp<="111";
	end if;
	if (ll=316 and cc>=138 and cc<148) then grbp<="111";
	end if;
	if (cc=187 and ll=316) then grbp<="111";
	end if;
	if (cc=197 and ll=316) then grbp<="111";
	end if;
	if (cc=200 and ll=316) then grbp<="111";
	end if;
	if (ll=316 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=221 and ll=316) then grbp<="111";
	end if;
	if (ll=316 and cc>=221 and cc<247) then grbp<="111";
	end if;
	if (cc=72 and ll=317) then grbp<="111";
	end if;
	if (cc=138 and ll=317) then grbp<="111";
	end if;
	if (ll=317 and cc>=138 and cc<148) then grbp<="111";
	end if;
	if (cc=197 and ll=317) then grbp<="111";
	end if;
	if (cc=199 and ll=317) then grbp<="111";
	end if;
	if (ll=317 and cc>=199 and cc<201) then grbp<="111";
	end if;
	if (cc=208 and ll=317) then grbp<="111";
	end if;
	if (cc=221 and ll=317) then grbp<="111";
	end if;
	if (ll=317 and cc>=221 and cc<245) then grbp<="111";
	end if;
	if (cc=26 and ll=318) then grbp<="111";
	end if;
	if (cc=67 and ll=318) then grbp<="111";
	end if;
	if (ll=318 and cc>=67 and cc<69) then grbp<="111";
	end if;
	if (cc=140 and ll=318) then grbp<="111";
	end if;
	if (ll=318 and cc>=140 and cc<145) then grbp<="111";
	end if;
	if (ll=318 and cc>=146 and cc<148) then grbp<="111";
	end if;
	if (cc=197 and ll=318) then grbp<="111";
	end if;
	if (cc=199 and ll=318) then grbp<="111";
	end if;
	if (cc=221 and ll=318) then grbp<="111";
	end if;
	if (ll=318 and cc>=221 and cc<244) then grbp<="111";
	end if;
	if (cc=56 and ll=319) then grbp<="111";
	end if;
	if (cc=72 and ll=319) then grbp<="111";
	end if;
	if (cc=140 and ll=319) then grbp<="111";
	end if;
	if (ll=319 and cc>=140 and cc<144) then grbp<="111";
	end if;
	if (cc=199 and ll=319) then grbp<="111";
	end if;
	if (cc=202 and ll=319) then grbp<="111";
	end if;
	if (cc=209 and ll=319) then grbp<="111";
	end if;
	if (cc=221 and ll=319) then grbp<="111";
	end if;
	if (ll=319 and cc>=221 and cc<242) then grbp<="111";
	end if;
	if (cc=35 and ll=320) then grbp<="111";
	end if;
	if (ll=320 and cc>=35 and cc<37) then grbp<="111";
	end if;
	if (cc=56 and ll=320) then grbp<="111";
	end if;
	if (ll=320 and cc>=56 and cc<58) then grbp<="111";
	end if;
	if (ll=320 and cc>=71 and cc<73) then grbp<="111";
	end if;
	if (ll=320 and cc>=75 and cc<77) then grbp<="111";
	end if;
	if (ll=320 and cc>=140 and cc<144) then grbp<="111";
	end if;
	if (cc=205 and ll=320) then grbp<="111";
	end if;
	if (ll=320 and cc>=205 and cc<208) then grbp<="111";
	end if;
	if (ll=320 and cc>=221 and cc<241) then grbp<="111";
	end if;
	if (cc=26 and ll=321) then grbp<="111";
	end if;
	if (cc=35 and ll=321) then grbp<="111";
	end if;
	if (cc=38 and ll=321) then grbp<="111";
	end if;
	if (cc=56 and ll=321) then grbp<="111";
	end if;
	if (cc=65 and ll=321) then grbp<="111";
	end if;
	if (cc=71 and ll=321) then grbp<="111";
	end if;
	if (ll=321 and cc>=71 and cc<73) then grbp<="111";
	end if;
	if (ll=321 and cc>=75 and cc<78) then grbp<="111";
	end if;
	if (cc=140 and ll=321) then grbp<="111";
	end if;
	if (ll=321 and cc>=140 and cc<147) then grbp<="111";
	end if;
	if (cc=205 and ll=321) then grbp<="111";
	end if;
	if (cc=220 and ll=321) then grbp<="111";
	end if;
	if (ll=321 and cc>=220 and cc<241) then grbp<="111";
	end if;
	if (cc=38 and ll=322) then grbp<="111";
	end if;
	if (cc=58 and ll=322) then grbp<="111";
	end if;
	if (cc=65 and ll=322) then grbp<="111";
	end if;
	if (cc=71 and ll=322) then grbp<="111";
	end if;
	if (ll=322 and cc>=71 and cc<73) then grbp<="111";
	end if;
	if (cc=136 and ll=322) then grbp<="111";
	end if;
	if (cc=138 and ll=322) then grbp<="111";
	end if;
	if (cc=140 and ll=322) then grbp<="111";
	end if;
	if (ll=322 and cc>=140 and cc<151) then grbp<="111";
	end if;
	if (cc=207 and ll=322) then grbp<="111";
	end if;
	if (cc=220 and ll=322) then grbp<="111";
	end if;
	if (ll=322 and cc>=220 and cc<239) then grbp<="111";
	end if;
	if (ll=323 and cc>=33 and cc<35) then grbp<="111";
	end if;
	if (cc=58 and ll=323) then grbp<="111";
	end if;
	if (cc=68 and ll=323) then grbp<="111";
	end if;
	if (cc=71 and ll=323) then grbp<="111";
	end if;
	if (ll=323 and cc>=71 and cc<73) then grbp<="111";
	end if;
	if (ll=323 and cc>=77 and cc<79) then grbp<="111";
	end if;
	if (ll=323 and cc>=143 and cc<153) then grbp<="111";
	end if;
	if (cc=207 and ll=323) then grbp<="111";
	end if;
	if (cc=220 and ll=323) then grbp<="111";
	end if;
	if (ll=323 and cc>=220 and cc<239) then grbp<="111";
	end if;
	if (cc=33 and ll=324) then grbp<="111";
	end if;
	if (cc=68 and ll=324) then grbp<="111";
	end if;
	if (cc=72 and ll=324) then grbp<="111";
	end if;
	if (ll=324 and cc>=72 and cc<74) then grbp<="111";
	end if;
	if (ll=324 and cc>=78 and cc<80) then grbp<="111";
	end if;
	if (cc=147 and ll=324) then grbp<="111";
	end if;
	if (ll=324 and cc>=147 and cc<155) then grbp<="111";
	end if;
	if (ll=324 and cc>=220 and cc<238) then grbp<="111";
	end if;
	if (ll=325 and cc>=32 and cc<34) then grbp<="111";
	end if;
	if (cc=67 and ll=325) then grbp<="111";
	end if;
	if (ll=325 and cc>=67 and cc<69) then grbp<="111";
	end if;
	if (cc=78 and ll=325) then grbp<="111";
	end if;
	if (ll=325 and cc>=78 and cc<80) then grbp<="111";
	end if;
	if (ll=325 and cc>=146 and cc<156) then grbp<="111";
	end if;
	if (ll=325 and cc>=220 and cc<239) then grbp<="111";
	end if;
	if (cc=31 and ll=326) then grbp<="111";
	end if;
	if (ll=326 and cc>=31 and cc<33) then grbp<="111";
	end if;
	if (cc=79 and ll=326) then grbp<="111";
	end if;
	if (ll=326 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=326 and cc>=146 and cc<157) then grbp<="111";
	end if;
	if (cc=220 and ll=326) then grbp<="111";
	end if;
	if (ll=326 and cc>=220 and cc<238) then grbp<="111";
	end if;
	if (cc=23 and ll=327) then grbp<="111";
	end if;
	if (cc=30 and ll=327) then grbp<="111";
	end if;
	if (ll=327 and cc>=30 and cc<32) then grbp<="111";
	end if;
	if (cc=67 and ll=327) then grbp<="111";
	end if;
	if (cc=80 and ll=327) then grbp<="111";
	end if;
	if (ll=327 and cc>=80 and cc<82) then grbp<="111";
	end if;
	if (ll=327 and cc>=146 and cc<159) then grbp<="111";
	end if;
	if (cc=220 and ll=327) then grbp<="111";
	end if;
	if (ll=327 and cc>=220 and cc<238) then grbp<="111";
	end if;
	if (ll=328 and cc>=29 and cc<31) then grbp<="111";
	end if;
	if (cc=61 and ll=328) then grbp<="111";
	end if;
	if (cc=66 and ll=328) then grbp<="111";
	end if;
	if (ll=328 and cc>=66 and cc<68) then grbp<="111";
	end if;
	if (cc=146 and ll=328) then grbp<="111";
	end if;
	if (ll=328 and cc>=146 and cc<160) then grbp<="111";
	end if;
	if (cc=220 and ll=328) then grbp<="111";
	end if;
	if (ll=328 and cc>=220 and cc<237) then grbp<="111";
	end if;
	if (ll=329 and cc>=28 and cc<31) then grbp<="111";
	end if;
	if (cc=78 and ll=329) then grbp<="111";
	end if;
	if (cc=82 and ll=329) then grbp<="111";
	end if;
	if (cc=146 and ll=329) then grbp<="111";
	end if;
	if (ll=329 and cc>=146 and cc<161) then grbp<="111";
	end if;
	if (cc=220 and ll=329) then grbp<="111";
	end if;
	if (ll=329 and cc>=220 and cc<236) then grbp<="111";
	end if;
	if (ll=330 and cc>=26 and cc<30) then grbp<="111";
	end if;
	if (cc=58 and ll=330) then grbp<="111";
	end if;
	if (cc=65 and ll=330) then grbp<="111";
	end if;
	if (ll=330 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (cc=82 and ll=330) then grbp<="111";
	end if;
	if (cc=146 and ll=330) then grbp<="111";
	end if;
	if (ll=330 and cc>=146 and cc<162) then grbp<="111";
	end if;
	if (cc=220 and ll=330) then grbp<="111";
	end if;
	if (ll=330 and cc>=220 and cc<235) then grbp<="111";
	end if;
	if (ll=331 and cc>=25 and cc<29) then grbp<="111";
	end if;
	if (cc=78 and ll=331) then grbp<="111";
	end if;
	if (cc=146 and ll=331) then grbp<="111";
	end if;
	if (ll=331 and cc>=146 and cc<163) then grbp<="111";
	end if;
	if (cc=221 and ll=331) then grbp<="111";
	end if;
	if (ll=331 and cc>=221 and cc<235) then grbp<="111";
	end if;
	if (cc=21 and ll=332) then grbp<="111";
	end if;
	if (cc=25 and ll=332) then grbp<="111";
	end if;
	if (ll=332 and cc>=25 and cc<28) then grbp<="111";
	end if;
	if (cc=78 and ll=332) then grbp<="111";
	end if;
	if (cc=83 and ll=332) then grbp<="111";
	end if;
	if (cc=146 and ll=332) then grbp<="111";
	end if;
	if (ll=332 and cc>=146 and cc<164) then grbp<="111";
	end if;
	if (cc=221 and ll=332) then grbp<="111";
	end if;
	if (ll=332 and cc>=221 and cc<235) then grbp<="111";
	end if;
	if (ll=333 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (cc=78 and ll=333) then grbp<="111";
	end if;
	if (cc=145 and ll=333) then grbp<="111";
	end if;
	if (ll=333 and cc>=145 and cc<165) then grbp<="111";
	end if;
	if (cc=220 and ll=333) then grbp<="111";
	end if;
	if (ll=333 and cc>=220 and cc<233) then grbp<="111";
	end if;
	if (cc=65 and ll=334) then grbp<="111";
	end if;
	if (cc=79 and ll=334) then grbp<="111";
	end if;
	if (cc=84 and ll=334) then grbp<="111";
	end if;
	if (cc=145 and ll=334) then grbp<="111";
	end if;
	if (ll=334 and cc>=145 and cc<166) then grbp<="111";
	end if;
	if (cc=220 and ll=334) then grbp<="111";
	end if;
	if (ll=334 and cc>=220 and cc<233) then grbp<="111";
	end if;
	if (cc=35 and ll=335) then grbp<="111";
	end if;
	if (cc=64 and ll=335) then grbp<="111";
	end if;
	if (cc=74 and ll=335) then grbp<="111";
	end if;
	if (cc=80 and ll=335) then grbp<="111";
	end if;
	if (cc=84 and ll=335) then grbp<="111";
	end if;
	if (cc=145 and ll=335) then grbp<="111";
	end if;
	if (ll=335 and cc>=145 and cc<167) then grbp<="111";
	end if;
	if (cc=220 and ll=335) then grbp<="111";
	end if;
	if (ll=335 and cc>=220 and cc<232) then grbp<="111";
	end if;
	if (cc=74 and ll=336) then grbp<="111";
	end if;
	if (cc=80 and ll=336) then grbp<="111";
	end if;
	if (cc=145 and ll=336) then grbp<="111";
	end if;
	if (ll=336 and cc>=145 and cc<168) then grbp<="111";
	end if;
	if (ll=336 and cc>=220 and cc<232) then grbp<="111";
	end if;
	if (cc=25 and ll=337) then grbp<="111";
	end if;
	if (cc=32 and ll=337) then grbp<="111";
	end if;
	if (cc=74 and ll=337) then grbp<="111";
	end if;
	if (ll=337 and cc>=74 and cc<76) then grbp<="111";
	end if;
	if (cc=145 and ll=337) then grbp<="111";
	end if;
	if (ll=337 and cc>=145 and cc<168) then grbp<="111";
	end if;
	if (ll=337 and cc>=220 and cc<231) then grbp<="111";
	end if;
	if (ll=338 and cc>=3 and cc<5) then grbp<="111";
	end if;
	if (cc=31 and ll=338) then grbp<="111";
	end if;
	if (ll=338 and cc>=31 and cc<33) then grbp<="111";
	end if;
	if (cc=74 and ll=338) then grbp<="111";
	end if;
	if (cc=81 and ll=338) then grbp<="111";
	end if;
	if (cc=85 and ll=338) then grbp<="111";
	end if;
	if (cc=144 and ll=338) then grbp<="111";
	end if;
	if (cc=146 and ll=338) then grbp<="111";
	end if;
	if (ll=338 and cc>=146 and cc<169) then grbp<="111";
	end if;
	if (ll=338 and cc>=220 and cc<231) then grbp<="111";
	end if;
	if (ll=339 and cc>=3 and cc<6) then grbp<="111";
	end if;
	if (ll=339 and cc>=31 and cc<33) then grbp<="111";
	end if;
	if (ll=339 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (cc=85 and ll=339) then grbp<="111";
	end if;
	if (cc=145 and ll=339) then grbp<="111";
	end if;
	if (ll=339 and cc>=145 and cc<170) then grbp<="111";
	end if;
	if (ll=339 and cc>=220 and cc<231) then grbp<="111";
	end if;
	if (ll=340 and cc>=2 and cc<7) then grbp<="111";
	end if;
	if (ll=340 and cc>=31 and cc<33) then grbp<="111";
	end if;
	if (ll=340 and cc>=76 and cc<79) then grbp<="111";
	end if;
	if (cc=146 and ll=340) then grbp<="111";
	end if;
	if (ll=340 and cc>=146 and cc<170) then grbp<="111";
	end if;
	if (cc=220 and ll=340) then grbp<="111";
	end if;
	if (ll=340 and cc>=220 and cc<231) then grbp<="111";
	end if;
	if (ll=341 and cc>=3 and cc<7) then grbp<="111";
	end if;
	if (ll=341 and cc>=31 and cc<33) then grbp<="111";
	end if;
	if (cc=78 and ll=341) then grbp<="111";
	end if;
	if (cc=82 and ll=341) then grbp<="111";
	end if;
	if (cc=86 and ll=341) then grbp<="111";
	end if;
	if (cc=144 and ll=341) then grbp<="111";
	end if;
	if (ll=341 and cc>=144 and cc<171) then grbp<="111";
	end if;
	if (cc=219 and ll=341) then grbp<="111";
	end if;
	if (ll=341 and cc>=219 and cc<230) then grbp<="111";
	end if;
	if (ll=342 and cc>=3 and cc<7) then grbp<="111";
	end if;
	if (cc=34 and ll=342) then grbp<="111";
	end if;
	if (cc=74 and ll=342) then grbp<="111";
	end if;
	if (cc=77 and ll=342) then grbp<="111";
	end if;
	if (cc=82 and ll=342) then grbp<="111";
	end if;
	if (ll=342 and cc>=82 and cc<84) then grbp<="111";
	end if;
	if (cc=145 and ll=342) then grbp<="111";
	end if;
	if (ll=342 and cc>=145 and cc<171) then grbp<="111";
	end if;
	if (ll=342 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=343 and cc>=3 and cc<9) then grbp<="111";
	end if;
	if (cc=34 and ll=343) then grbp<="111";
	end if;
	if (cc=83 and ll=343) then grbp<="111";
	end if;
	if (cc=86 and ll=343) then grbp<="111";
	end if;
	if (cc=146 and ll=343) then grbp<="111";
	end if;
	if (ll=343 and cc>=146 and cc<172) then grbp<="111";
	end if;
	if (ll=343 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=344 and cc>=4 and cc<9) then grbp<="111";
	end if;
	if (cc=31 and ll=344) then grbp<="111";
	end if;
	if (cc=34 and ll=344) then grbp<="111";
	end if;
	if (cc=86 and ll=344) then grbp<="111";
	end if;
	if (cc=147 and ll=344) then grbp<="111";
	end if;
	if (ll=344 and cc>=147 and cc<172) then grbp<="111";
	end if;
	if (cc=219 and ll=344) then grbp<="111";
	end if;
	if (ll=344 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=345 and cc>=4 and cc<9) then grbp<="111";
	end if;
	if (cc=74 and ll=345) then grbp<="111";
	end if;
	if (cc=84 and ll=345) then grbp<="111";
	end if;
	if (cc=87 and ll=345) then grbp<="111";
	end if;
	if (cc=148 and ll=345) then grbp<="111";
	end if;
	if (ll=345 and cc>=148 and cc<173) then grbp<="111";
	end if;
	if (cc=219 and ll=345) then grbp<="111";
	end if;
	if (ll=345 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=346 and cc>=5 and cc<10) then grbp<="111";
	end if;
	if (cc=31 and ll=346) then grbp<="111";
	end if;
	if (cc=79 and ll=346) then grbp<="111";
	end if;
	if (cc=84 and ll=346) then grbp<="111";
	end if;
	if (cc=87 and ll=346) then grbp<="111";
	end if;
	if (cc=149 and ll=346) then grbp<="111";
	end if;
	if (ll=346 and cc>=149 and cc<173) then grbp<="111";
	end if;
	if (cc=219 and ll=346) then grbp<="111";
	end if;
	if (ll=346 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=347 and cc>=5 and cc<10) then grbp<="111";
	end if;
	if (ll=347 and cc>=20 and cc<22) then grbp<="111";
	end if;
	if (cc=79 and ll=347) then grbp<="111";
	end if;
	if (ll=347 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=87 and ll=347) then grbp<="111";
	end if;
	if (cc=149 and ll=347) then grbp<="111";
	end if;
	if (ll=347 and cc>=149 and cc<173) then grbp<="111";
	end if;
	if (cc=219 and ll=347) then grbp<="111";
	end if;
	if (ll=347 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=348 and cc>=5 and cc<10) then grbp<="111";
	end if;
	if (cc=79 and ll=348) then grbp<="111";
	end if;
	if (ll=348 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=149 and ll=348) then grbp<="111";
	end if;
	if (ll=348 and cc>=149 and cc<174) then grbp<="111";
	end if;
	if (ll=348 and cc>=219 and cc<229) then grbp<="111";
	end if;
	if (ll=349 and cc>=5 and cc<10) then grbp<="111";
	end if;
	if (cc=79 and ll=349) then grbp<="111";
	end if;
	if (ll=349 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=149 and ll=349) then grbp<="111";
	end if;
	if (ll=349 and cc>=149 and cc<174) then grbp<="111";
	end if;
	if (ll=349 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=350 and cc>=5 and cc<10) then grbp<="111";
	end if;
	if (cc=22 and ll=350) then grbp<="111";
	end if;
	if (cc=24 and ll=350) then grbp<="111";
	end if;
	if (cc=79 and ll=350) then grbp<="111";
	end if;
	if (ll=350 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=147 and ll=350) then grbp<="111";
	end if;
	if (cc=150 and ll=350) then grbp<="111";
	end if;
	if (ll=350 and cc>=150 and cc<174) then grbp<="111";
	end if;
	if (ll=350 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=351 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=79 and ll=351) then grbp<="111";
	end if;
	if (ll=351 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=148 and ll=351) then grbp<="111";
	end if;
	if (cc=150 and ll=351) then grbp<="111";
	end if;
	if (ll=351 and cc>=150 and cc<175) then grbp<="111";
	end if;
	if (ll=351 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (ll=352 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=76 and ll=352) then grbp<="111";
	end if;
	if (cc=78 and ll=352) then grbp<="111";
	end if;
	if (cc=80 and ll=352) then grbp<="111";
	end if;
	if (cc=87 and ll=352) then grbp<="111";
	end if;
	if (cc=149 and ll=352) then grbp<="111";
	end if;
	if (ll=352 and cc>=149 and cc<175) then grbp<="111";
	end if;
	if (ll=352 and cc>=217 and cc<227) then grbp<="111";
	end if;
	if (ll=353 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (ll=353 and cc>=77 and cc<80) then grbp<="111";
	end if;
	if (ll=353 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (ll=353 and cc>=149 and cc<175) then grbp<="111";
	end if;
	if (ll=353 and cc>=215 and cc<227) then grbp<="111";
	end if;
	if (ll=354 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=77 and ll=354) then grbp<="111";
	end if;
	if (ll=354 and cc>=77 and cc<81) then grbp<="111";
	end if;
	if (ll=354 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (ll=354 and cc>=150 and cc<176) then grbp<="111";
	end if;
	if (ll=354 and cc>=215 and cc<227) then grbp<="111";
	end if;
	if (ll=355 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=23 and ll=355) then grbp<="111";
	end if;
	if (cc=33 and ll=355) then grbp<="111";
	end if;
	if (cc=51 and ll=355) then grbp<="111";
	end if;
	if (cc=77 and ll=355) then grbp<="111";
	end if;
	if (ll=355 and cc>=77 and cc<79) then grbp<="111";
	end if;
	if (cc=86 and ll=355) then grbp<="111";
	end if;
	if (ll=355 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (cc=151 and ll=355) then grbp<="111";
	end if;
	if (ll=355 and cc>=151 and cc<176) then grbp<="111";
	end if;
	if (ll=355 and cc>=214 and cc<226) then grbp<="111";
	end if;
	if (ll=356 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=77 and ll=356) then grbp<="111";
	end if;
	if (cc=80 and ll=356) then grbp<="111";
	end if;
	if (cc=86 and ll=356) then grbp<="111";
	end if;
	if (ll=356 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (ll=356 and cc>=150 and cc<176) then grbp<="111";
	end if;
	if (ll=356 and cc>=213 and cc<226) then grbp<="111";
	end if;
	if (ll=357 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=86 and ll=357) then grbp<="111";
	end if;
	if (ll=357 and cc>=86 and cc<88) then grbp<="111";
	end if;
	if (cc=151 and ll=357) then grbp<="111";
	end if;
	if (ll=357 and cc>=151 and cc<176) then grbp<="111";
	end if;
	if (ll=357 and cc>=212 and cc<226) then grbp<="111";
	end if;
	if (ll=358 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (ll=358 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=149 and ll=358) then grbp<="111";
	end if;
	if (ll=358 and cc>=149 and cc<177) then grbp<="111";
	end if;
	if (ll=358 and cc>=212 and cc<225) then grbp<="111";
	end if;
	if (ll=359 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (ll=359 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (cc=86 and ll=359) then grbp<="111";
	end if;
	if (cc=88 and ll=359) then grbp<="111";
	end if;
	if (cc=150 and ll=359) then grbp<="111";
	end if;
	if (ll=359 and cc>=150 and cc<177) then grbp<="111";
	end if;
	if (ll=359 and cc>=211 and cc<225) then grbp<="111";
	end if;
	if (ll=360 and cc>=5 and cc<11) then grbp<="111";
	end if;
	if (cc=79 and ll=360) then grbp<="111";
	end if;
	if (cc=82 and ll=360) then grbp<="111";
	end if;
	if (cc=85 and ll=360) then grbp<="111";
	end if;
	if (ll=360 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (cc=152 and ll=360) then grbp<="111";
	end if;
	if (ll=360 and cc>=152 and cc<177) then grbp<="111";
	end if;
	if (ll=360 and cc>=211 and cc<225) then grbp<="111";
	end if;
	if (ll=361 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=79 and ll=361) then grbp<="111";
	end if;
	if (cc=85 and ll=361) then grbp<="111";
	end if;
	if (ll=361 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (cc=150 and ll=361) then grbp<="111";
	end if;
	if (ll=361 and cc>=150 and cc<152) then grbp<="111";
	end if;
	if (ll=361 and cc>=153 and cc<177) then grbp<="111";
	end if;
	if (cc=211 and ll=361) then grbp<="111";
	end if;
	if (ll=361 and cc>=211 and cc<224) then grbp<="111";
	end if;
	if (ll=362 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=78 and ll=362) then grbp<="111";
	end if;
	if (ll=362 and cc>=78 and cc<81) then grbp<="111";
	end if;
	if (ll=362 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (cc=152 and ll=362) then grbp<="111";
	end if;
	if (ll=362 and cc>=152 and cc<177) then grbp<="111";
	end if;
	if (ll=362 and cc>=211 and cc<224) then grbp<="111";
	end if;
	if (ll=363 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=78 and ll=363) then grbp<="111";
	end if;
	if (ll=363 and cc>=78 and cc<81) then grbp<="111";
	end if;
	if (ll=363 and cc>=84 and cc<86) then grbp<="111";
	end if;
	if (ll=363 and cc>=151 and cc<178) then grbp<="111";
	end if;
	if (ll=363 and cc>=211 and cc<224) then grbp<="111";
	end if;
	if (ll=364 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=82 and ll=364) then grbp<="111";
	end if;
	if (ll=364 and cc>=82 and cc<86) then grbp<="111";
	end if;
	if (ll=364 and cc>=151 and cc<178) then grbp<="111";
	end if;
	if (ll=364 and cc>=211 and cc<224) then grbp<="111";
	end if;
	if (ll=365 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=83 and ll=365) then grbp<="111";
	end if;
	if (ll=365 and cc>=83 and cc<86) then grbp<="111";
	end if;
	if (ll=365 and cc>=151 and cc<178) then grbp<="111";
	end if;
	if (ll=365 and cc>=211 and cc<223) then grbp<="111";
	end if;
	if (ll=366 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (ll=366 and cc>=83 and cc<87) then grbp<="111";
	end if;
	if (ll=366 and cc>=152 and cc<178) then grbp<="111";
	end if;
	if (ll=366 and cc>=210 and cc<223) then grbp<="111";
	end if;
	if (ll=367 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=83 and ll=367) then grbp<="111";
	end if;
	if (cc=85 and ll=367) then grbp<="111";
	end if;
	if (ll=367 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (cc=153 and ll=367) then grbp<="111";
	end if;
	if (ll=367 and cc>=153 and cc<178) then grbp<="111";
	end if;
	if (ll=367 and cc>=211 and cc<223) then grbp<="111";
	end if;
	if (ll=368 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (ll=368 and cc>=21 and cc<27) then grbp<="111";
	end if;
	if (cc=153 and ll=368) then grbp<="111";
	end if;
	if (ll=368 and cc>=153 and cc<178) then grbp<="111";
	end if;
	if (ll=368 and cc>=211 and cc<223) then grbp<="111";
	end if;
	if (ll=369 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (ll=369 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (ll=369 and cc>=152 and cc<179) then grbp<="111";
	end if;
	if (ll=369 and cc>=210 and cc<222) then grbp<="111";
	end if;
	if (ll=370 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=94 and ll=370) then grbp<="111";
	end if;
	if (cc=153 and ll=370) then grbp<="111";
	end if;
	if (ll=370 and cc>=153 and cc<179) then grbp<="111";
	end if;
	if (ll=370 and cc>=210 and cc<222) then grbp<="111";
	end if;
	if (ll=371 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (ll=371 and cc>=154 and cc<179) then grbp<="111";
	end if;
	if (cc=210 and ll=371) then grbp<="111";
	end if;
	if (ll=371 and cc>=210 and cc<222) then grbp<="111";
	end if;
	if (ll=372 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=31 and ll=372) then grbp<="111";
	end if;
	if (cc=154 and ll=372) then grbp<="111";
	end if;
	if (ll=372 and cc>=154 and cc<179) then grbp<="111";
	end if;
	if (cc=211 and ll=372) then grbp<="111";
	end if;
	if (ll=372 and cc>=211 and cc<222) then grbp<="111";
	end if;
	if (ll=373 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=152 and ll=373) then grbp<="111";
	end if;
	if (cc=154 and ll=373) then grbp<="111";
	end if;
	if (ll=373 and cc>=154 and cc<179) then grbp<="111";
	end if;
	if (ll=373 and cc>=211 and cc<221) then grbp<="111";
	end if;
	if (ll=374 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=81 and ll=374) then grbp<="111";
	end if;
	if (cc=151 and ll=374) then grbp<="111";
	end if;
	if (ll=374 and cc>=151 and cc<153) then grbp<="111";
	end if;
	if (ll=374 and cc>=155 and cc<179) then grbp<="111";
	end if;
	if (cc=214 and ll=374) then grbp<="111";
	end if;
	if (ll=374 and cc>=214 and cc<221) then grbp<="111";
	end if;
	if (ll=375 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=76 and ll=375) then grbp<="111";
	end if;
	if (cc=82 and ll=375) then grbp<="111";
	end if;
	if (cc=152 and ll=375) then grbp<="111";
	end if;
	if (ll=375 and cc>=152 and cc<180) then grbp<="111";
	end if;
	if (ll=375 and cc>=216 and cc<221) then grbp<="111";
	end if;
	if (ll=376 and cc>=6 and cc<12) then grbp<="111";
	end if;
	if (cc=31 and ll=376) then grbp<="111";
	end if;
	if (cc=153 and ll=376) then grbp<="111";
	end if;
	if (cc=156 and ll=376) then grbp<="111";
	end if;
	if (ll=376 and cc>=156 and cc<180) then grbp<="111";
	end if;
	if (ll=376 and cc>=216 and cc<221) then grbp<="111";
	end if;
	if (ll=377 and cc>=6 and cc<11) then grbp<="111";
	end if;
	if (cc=73 and ll=377) then grbp<="111";
	end if;
	if (ll=377 and cc>=73 and cc<75) then grbp<="111";
	end if;
	if (ll=377 and cc>=156 and cc<180) then grbp<="111";
	end if;
	if (ll=377 and cc>=215 and cc<221) then grbp<="111";
	end if;
	if (ll=378 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=86 and ll=378) then grbp<="111";
	end if;
	if (cc=156 and ll=378) then grbp<="111";
	end if;
	if (ll=378 and cc>=156 and cc<180) then grbp<="111";
	end if;
	if (ll=378 and cc>=215 and cc<221) then grbp<="111";
	end if;
	if (ll=379 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=86 and ll=379) then grbp<="111";
	end if;
	if (cc=156 and ll=379) then grbp<="111";
	end if;
	if (ll=379 and cc>=156 and cc<180) then grbp<="111";
	end if;
	if (ll=379 and cc>=215 and cc<221) then grbp<="111";
	end if;
	if (ll=380 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (ll=380 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (cc=84 and ll=380) then grbp<="111";
	end if;
	if (ll=380 and cc>=84 and cc<86) then grbp<="111";
	end if;
	if (ll=380 and cc>=156 and cc<181) then grbp<="111";
	end if;
	if (ll=380 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=381 and cc>=6 and cc<12) then grbp<="111";
	end if;
	if (cc=84 and ll=381) then grbp<="111";
	end if;
	if (ll=381 and cc>=84 and cc<86) then grbp<="111";
	end if;
	if (ll=381 and cc>=154 and cc<181) then grbp<="111";
	end if;
	if (cc=215 and ll=381) then grbp<="111";
	end if;
	if (ll=381 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=382 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=157 and ll=382) then grbp<="111";
	end if;
	if (ll=382 and cc>=157 and cc<181) then grbp<="111";
	end if;
	if (ll=382 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=383 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (ll=383 and cc>=158 and cc<181) then grbp<="111";
	end if;
	if (ll=383 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=384 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (ll=384 and cc>=158 and cc<181) then grbp<="111";
	end if;
	if (ll=384 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=385 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=159 and ll=385) then grbp<="111";
	end if;
	if (ll=385 and cc>=159 and cc<181) then grbp<="111";
	end if;
	if (ll=385 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=386 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=72 and ll=386) then grbp<="111";
	end if;
	if (cc=158 and ll=386) then grbp<="111";
	end if;
	if (ll=386 and cc>=158 and cc<182) then grbp<="111";
	end if;
	if (ll=386 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=387 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=156 and ll=387) then grbp<="111";
	end if;
	if (ll=387 and cc>=156 and cc<158) then grbp<="111";
	end if;
	if (ll=387 and cc>=159 and cc<182) then grbp<="111";
	end if;
	if (ll=387 and cc>=214 and cc<218) then grbp<="111";
	end if;
	if (ll=388 and cc>=7 and cc<12) then grbp<="111";
	end if;
	if (cc=159 and ll=388) then grbp<="111";
	end if;
	if (ll=388 and cc>=159 and cc<182) then grbp<="111";
	end if;
	if (ll=388 and cc>=214 and cc<218) then grbp<="111";
	end if;
	if (ll=389 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=160 and ll=389) then grbp<="111";
	end if;
	if (ll=389 and cc>=160 and cc<182) then grbp<="111";
	end if;
	if (ll=389 and cc>=214 and cc<218) then grbp<="111";
	end if;
	if (ll=390 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=74 and ll=390) then grbp<="111";
	end if;
	if (cc=159 and ll=390) then grbp<="111";
	end if;
	if (ll=390 and cc>=159 and cc<182) then grbp<="111";
	end if;
	if (ll=390 and cc>=213 and cc<218) then grbp<="111";
	end if;
	if (ll=391 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=159 and ll=391) then grbp<="111";
	end if;
	if (ll=391 and cc>=159 and cc<182) then grbp<="111";
	end if;
	if (ll=391 and cc>=213 and cc<218) then grbp<="111";
	end if;
	if (ll=392 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=160 and ll=392) then grbp<="111";
	end if;
	if (ll=392 and cc>=160 and cc<183) then grbp<="111";
	end if;
	if (cc=213 and ll=392) then grbp<="111";
	end if;
	if (ll=392 and cc>=213 and cc<217) then grbp<="111";
	end if;
	if (ll=393 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=393 and cc>=73 and cc<75) then grbp<="111";
	end if;
	if (ll=393 and cc>=160 and cc<183) then grbp<="111";
	end if;
	if (ll=393 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=393 and cc>=213 and cc<217) then grbp<="111";
	end if;
	if (ll=394 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=160 and ll=394) then grbp<="111";
	end if;
	if (ll=394 and cc>=160 and cc<183) then grbp<="111";
	end if;
	if (ll=394 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=394 and cc>=213 and cc<217) then grbp<="111";
	end if;
	if (ll=395 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=161 and ll=395) then grbp<="111";
	end if;
	if (cc=163 and ll=395) then grbp<="111";
	end if;
	if (ll=395 and cc>=163 and cc<183) then grbp<="111";
	end if;
	if (ll=395 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=395 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (ll=396 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=76 and ll=396) then grbp<="111";
	end if;
	if (cc=160 and ll=396) then grbp<="111";
	end if;
	if (ll=396 and cc>=160 and cc<183) then grbp<="111";
	end if;
	if (ll=396 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=396 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (ll=397 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=397 and cc>=76 and cc<78) then grbp<="111";
	end if;
	if (ll=397 and cc>=160 and cc<183) then grbp<="111";
	end if;
	if (ll=397 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=398 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=398 and cc>=162 and cc<184) then grbp<="111";
	end if;
	if (cc=7 and ll=399) then grbp<="111";
	end if;
	if (ll=399 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=399 and cc>=162 and cc<184) then grbp<="111";
	end if;
	if (ll=399 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=400 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=400 and cc>=159 and cc<161) then grbp<="111";
	end if;
	if (ll=400 and cc>=163 and cc<184) then grbp<="111";
	end if;
	if (ll=400 and cc>=207 and cc<211) then grbp<="111";
	end if;
	if (ll=401 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=162 and ll=401) then grbp<="111";
	end if;
	if (ll=401 and cc>=162 and cc<184) then grbp<="111";
	end if;
	if (ll=401 and cc>=207 and cc<211) then grbp<="111";
	end if;
	if (ll=402 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (ll=402 and cc>=162 and cc<184) then grbp<="111";
	end if;
	if (ll=402 and cc>=207 and cc<211) then grbp<="111";
	end if;
	if (ll=403 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=76 and ll=403) then grbp<="111";
	end if;
	if (cc=151 and ll=403) then grbp<="111";
	end if;
	if (cc=153 and ll=403) then grbp<="111";
	end if;
	if (cc=158 and ll=403) then grbp<="111";
	end if;
	if (cc=162 and ll=403) then grbp<="111";
	end if;
	if (ll=403 and cc>=162 and cc<184) then grbp<="111";
	end if;
	if (ll=403 and cc>=207 and cc<211) then grbp<="111";
	end if;
	if (ll=404 and cc>=7 and cc<13) then grbp<="111";
	end if;
	if (cc=136 and ll=404) then grbp<="111";
	end if;
	if (cc=138 and ll=404) then grbp<="111";
	end if;
	if (cc=151 and ll=404) then grbp<="111";
	end if;
	if (cc=153 and ll=404) then grbp<="111";
	end if;
	if (ll=404 and cc>=153 and cc<155) then grbp<="111";
	end if;
	if (cc=162 and ll=404) then grbp<="111";
	end if;
	if (ll=404 and cc>=162 and cc<185) then grbp<="111";
	end if;
	if (ll=404 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (cc=221 and ll=404) then grbp<="111";
	end if;
	if (ll=404 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=404 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=404 and cc>=234 and cc<236) then grbp<="111";
	end if;
	if (ll=404 and cc>=238 and cc<241) then grbp<="111";
	end if;
	if (ll=404 and cc>=243 and cc<245) then grbp<="111";
	end if;
	if (ll=405 and cc>=8 and cc<13) then grbp<="111";
	end if;
	if (cc=26 and ll=405) then grbp<="111";
	end if;
	if (cc=131 and ll=405) then grbp<="111";
	end if;
	if (cc=136 and ll=405) then grbp<="111";
	end if;
	if (cc=138 and ll=405) then grbp<="111";
	end if;
	if (cc=151 and ll=405) then grbp<="111";
	end if;
	if (cc=153 and ll=405) then grbp<="111";
	end if;
	if (ll=405 and cc>=153 and cc<155) then grbp<="111";
	end if;
	if (cc=160 and ll=405) then grbp<="111";
	end if;
	if (cc=163 and ll=405) then grbp<="111";
	end if;
	if (ll=405 and cc>=163 and cc<185) then grbp<="111";
	end if;
	if (cc=207 and ll=405) then grbp<="111";
	end if;
	if (ll=405 and cc>=207 and cc<211) then grbp<="111";
	end if;
	if (cc=217 and ll=405) then grbp<="111";
	end if;
	if (cc=220 and ll=405) then grbp<="111";
	end if;
	if (cc=222 and ll=405) then grbp<="111";
	end if;
	if (cc=225 and ll=405) then grbp<="111";
	end if;
	if (cc=227 and ll=405) then grbp<="111";
	end if;
	if (cc=230 and ll=405) then grbp<="111";
	end if;
	if (cc=234 and ll=405) then grbp<="111";
	end if;
	if (cc=236 and ll=405) then grbp<="111";
	end if;
	if (cc=238 and ll=405) then grbp<="111";
	end if;
	if (cc=240 and ll=405) then grbp<="111";
	end if;
	if (cc=242 and ll=405) then grbp<="111";
	end if;
	if (cc=8 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=8 and cc<13) then grbp<="111";
	end if;
	if (cc=77 and ll=406) then grbp<="111";
	end if;
	if (cc=131 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=131 and cc<134) then grbp<="111";
	end if;
	if (ll=406 and cc>=135 and cc<139) then grbp<="111";
	end if;
	if (ll=406 and cc>=141 and cc<143) then grbp<="111";
	end if;
	if (ll=406 and cc>=145 and cc<147) then grbp<="111";
	end if;
	if (cc=152 and ll=406) then grbp<="111";
	end if;
	if (cc=154 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=154 and cc<157) then grbp<="111";
	end if;
	if (cc=160 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=160 and cc<186) then grbp<="111";
	end if;
	if (cc=195 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=195 and cc<197) then grbp<="111";
	end if;
	if (ll=406 and cc>=198 and cc<200) then grbp<="111";
	end if;
	if (cc=207 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=406 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=220 and ll=406) then grbp<="111";
	end if;
	if (cc=227 and ll=406) then grbp<="111";
	end if;
	if (cc=229 and ll=406) then grbp<="111";
	end if;
	if (ll=406 and cc>=229 and cc<231) then grbp<="111";
	end if;
	if (cc=236 and ll=406) then grbp<="111";
	end if;
	if (cc=240 and ll=406) then grbp<="111";
	end if;
	if (cc=242 and ll=406) then grbp<="111";
	end if;
	if (cc=245 and ll=406) then grbp<="111";
	end if;
	if (cc=8 and ll=407) then grbp<="111";
	end if;
	if (ll=407 and cc>=8 and cc<13) then grbp<="111";
	end if;
	if (ll=407 and cc>=77 and cc<79) then grbp<="111";
	end if;
	if (ll=407 and cc>=131 and cc<139) then grbp<="111";
	end if;
	if (ll=407 and cc>=140 and cc<143) then grbp<="111";
	end if;
	if (ll=407 and cc>=144 and cc<147) then grbp<="111";
	end if;
	if (cc=150 and ll=407) then grbp<="111";
	end if;
	if (cc=152 and ll=407) then grbp<="111";
	end if;
	if (cc=154 and ll=407) then grbp<="111";
	end if;
	if (ll=407 and cc>=154 and cc<157) then grbp<="111";
	end if;
	if (cc=160 and ll=407) then grbp<="111";
	end if;
	if (ll=407 and cc>=160 and cc<186) then grbp<="111";
	end if;
	if (cc=192 and ll=407) then grbp<="111";
	end if;
	if (cc=194 and ll=407) then grbp<="111";
	end if;
	if (ll=407 and cc>=194 and cc<197) then grbp<="111";
	end if;
	if (ll=407 and cc>=198 and cc<200) then grbp<="111";
	end if;
	if (ll=407 and cc>=201 and cc<203) then grbp<="111";
	end if;
	if (cc=207 and ll=407) then grbp<="111";
	end if;
	if (cc=209 and ll=407) then grbp<="111";
	end if;
	if (cc=213 and ll=407) then grbp<="111";
	end if;
	if (cc=220 and ll=407) then grbp<="111";
	end if;
	if (cc=223 and ll=407) then grbp<="111";
	end if;
	if (ll=407 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=233 and ll=407) then grbp<="111";
	end if;
	if (cc=240 and ll=407) then grbp<="111";
	end if;
	if (cc=242 and ll=407) then grbp<="111";
	end if;
	if (cc=245 and ll=407) then grbp<="111";
	end if;
	if (cc=8 and ll=408) then grbp<="111";
	end if;
	if (ll=408 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (cc=131 and ll=408) then grbp<="111";
	end if;
	if (cc=134 and ll=408) then grbp<="111";
	end if;
	if (cc=136 and ll=408) then grbp<="111";
	end if;
	if (cc=138 and ll=408) then grbp<="111";
	end if;
	if (cc=140 and ll=408) then grbp<="111";
	end if;
	if (cc=142 and ll=408) then grbp<="111";
	end if;
	if (cc=144 and ll=408) then grbp<="111";
	end if;
	if (cc=150 and ll=408) then grbp<="111";
	end if;
	if (cc=152 and ll=408) then grbp<="111";
	end if;
	if (cc=154 and ll=408) then grbp<="111";
	end if;
	if (cc=156 and ll=408) then grbp<="111";
	end if;
	if (ll=408 and cc>=156 and cc<159) then grbp<="111";
	end if;
	if (cc=163 and ll=408) then grbp<="111";
	end if;
	if (ll=408 and cc>=163 and cc<185) then grbp<="111";
	end if;
	if (cc=190 and ll=408) then grbp<="111";
	end if;
	if (cc=192 and ll=408) then grbp<="111";
	end if;
	if (cc=194 and ll=408) then grbp<="111";
	end if;
	if (cc=197 and ll=408) then grbp<="111";
	end if;
	if (cc=202 and ll=408) then grbp<="111";
	end if;
	if (cc=205 and ll=408) then grbp<="111";
	end if;
	if (cc=207 and ll=408) then grbp<="111";
	end if;
	if (cc=213 and ll=408) then grbp<="111";
	end if;
	if (cc=216 and ll=408) then grbp<="111";
	end if;
	if (cc=220 and ll=408) then grbp<="111";
	end if;
	if (cc=223 and ll=408) then grbp<="111";
	end if;
	if (ll=408 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (ll=408 and cc>=233 and cc<237) then grbp<="111";
	end if;
	if (ll=408 and cc>=239 and cc<241) then grbp<="111";
	end if;
	if (cc=245 and ll=408) then grbp<="111";
	end if;
	if (cc=8 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (cc=26 and ll=409) then grbp<="111";
	end if;
	if (cc=131 and ll=409) then grbp<="111";
	end if;
	if (cc=134 and ll=409) then grbp<="111";
	end if;
	if (cc=136 and ll=409) then grbp<="111";
	end if;
	if (cc=138 and ll=409) then grbp<="111";
	end if;
	if (cc=142 and ll=409) then grbp<="111";
	end if;
	if (cc=144 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=144 and cc<147) then grbp<="111";
	end if;
	if (cc=152 and ll=409) then grbp<="111";
	end if;
	if (cc=154 and ll=409) then grbp<="111";
	end if;
	if (cc=156 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=156 and cc<159) then grbp<="111";
	end if;
	if (cc=163 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=163 and cc<185) then grbp<="111";
	end if;
	if (cc=192 and ll=409) then grbp<="111";
	end if;
	if (cc=194 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=194 and cc<198) then grbp<="111";
	end if;
	if (cc=202 and ll=409) then grbp<="111";
	end if;
	if (cc=205 and ll=409) then grbp<="111";
	end if;
	if (cc=213 and ll=409) then grbp<="111";
	end if;
	if (cc=220 and ll=409) then grbp<="111";
	end if;
	if (cc=223 and ll=409) then grbp<="111";
	end if;
	if (ll=409 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=233 and ll=409) then grbp<="111";
	end if;
	if (cc=236 and ll=409) then grbp<="111";
	end if;
	if (cc=240 and ll=409) then grbp<="111";
	end if;
	if (cc=242 and ll=409) then grbp<="111";
	end if;
	if (cc=245 and ll=409) then grbp<="111";
	end if;
	if (cc=8 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (cc=26 and ll=410) then grbp<="111";
	end if;
	if (cc=131 and ll=410) then grbp<="111";
	end if;
	if (cc=134 and ll=410) then grbp<="111";
	end if;
	if (cc=136 and ll=410) then grbp<="111";
	end if;
	if (cc=138 and ll=410) then grbp<="111";
	end if;
	if (cc=142 and ll=410) then grbp<="111";
	end if;
	if (cc=145 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=145 and cc<147) then grbp<="111";
	end if;
	if (cc=152 and ll=410) then grbp<="111";
	end if;
	if (cc=154 and ll=410) then grbp<="111";
	end if;
	if (cc=157 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=157 and cc<159) then grbp<="111";
	end if;
	if (cc=162 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=162 and cc<187) then grbp<="111";
	end if;
	if (cc=194 and ll=410) then grbp<="111";
	end if;
	if (cc=199 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=199 and cc<201) then grbp<="111";
	end if;
	if (cc=205 and ll=410) then grbp<="111";
	end if;
	if (cc=207 and ll=410) then grbp<="111";
	end if;
	if (cc=213 and ll=410) then grbp<="111";
	end if;
	if (cc=215 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=215 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=410) then grbp<="111";
	end if;
	if (ll=410 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=233 and ll=410) then grbp<="111";
	end if;
	if (cc=236 and ll=410) then grbp<="111";
	end if;
	if (cc=242 and ll=410) then grbp<="111";
	end if;
	if (cc=245 and ll=410) then grbp<="111";
	end if;
	if (cc=8 and ll=411) then grbp<="111";
	end if;
	if (ll=411 and cc>=8 and cc<13) then grbp<="111";
	end if;
	if (cc=131 and ll=411) then grbp<="111";
	end if;
	if (cc=134 and ll=411) then grbp<="111";
	end if;
	if (cc=136 and ll=411) then grbp<="111";
	end if;
	if (cc=138 and ll=411) then grbp<="111";
	end if;
	if (cc=140 and ll=411) then grbp<="111";
	end if;
	if (cc=142 and ll=411) then grbp<="111";
	end if;
	if (cc=144 and ll=411) then grbp<="111";
	end if;
	if (cc=146 and ll=411) then grbp<="111";
	end if;
	if (cc=150 and ll=411) then grbp<="111";
	end if;
	if (cc=154 and ll=411) then grbp<="111";
	end if;
	if (cc=156 and ll=411) then grbp<="111";
	end if;
	if (cc=158 and ll=411) then grbp<="111";
	end if;
	if (cc=160 and ll=411) then grbp<="111";
	end if;
	if (cc=162 and ll=411) then grbp<="111";
	end if;
	if (ll=411 and cc>=162 and cc<187) then grbp<="111";
	end if;
	if (cc=194 and ll=411) then grbp<="111";
	end if;
	if (cc=197 and ll=411) then grbp<="111";
	end if;
	if (cc=199 and ll=411) then grbp<="111";
	end if;
	if (ll=411 and cc>=199 and cc<201) then grbp<="111";
	end if;
	if (cc=205 and ll=411) then grbp<="111";
	end if;
	if (cc=207 and ll=411) then grbp<="111";
	end if;
	if (cc=209 and ll=411) then grbp<="111";
	end if;
	if (cc=213 and ll=411) then grbp<="111";
	end if;
	if (cc=218 and ll=411) then grbp<="111";
	end if;
	if (cc=220 and ll=411) then grbp<="111";
	end if;
	if (cc=223 and ll=411) then grbp<="111";
	end if;
	if (ll=411 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=233 and ll=411) then grbp<="111";
	end if;
	if (cc=236 and ll=411) then grbp<="111";
	end if;
	if (cc=240 and ll=411) then grbp<="111";
	end if;
	if (cc=242 and ll=411) then grbp<="111";
	end if;
	if (cc=8 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (ll=412 and cc>=22 and cc<25) then grbp<="111";
	end if;
	if (cc=131 and ll=412) then grbp<="111";
	end if;
	if (cc=134 and ll=412) then grbp<="111";
	end if;
	if (cc=136 and ll=412) then grbp<="111";
	end if;
	if (cc=138 and ll=412) then grbp<="111";
	end if;
	if (cc=140 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=140 and cc<143) then grbp<="111";
	end if;
	if (ll=412 and cc>=144 and cc<147) then grbp<="111";
	end if;
	if (ll=412 and cc>=148 and cc<150) then grbp<="111";
	end if;
	if (cc=154 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=154 and cc<157) then grbp<="111";
	end if;
	if (cc=160 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=160 and cc<187) then grbp<="111";
	end if;
	if (cc=192 and ll=412) then grbp<="111";
	end if;
	if (cc=194 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=194 and cc<197) then grbp<="111";
	end if;
	if (ll=412 and cc>=199 and cc<201) then grbp<="111";
	end if;
	if (ll=412 and cc>=203 and cc<206) then grbp<="111";
	end if;
	if (ll=412 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (cc=221 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (cc=227 and ll=412) then grbp<="111";
	end if;
	if (cc=234 and ll=412) then grbp<="111";
	end if;
	if (ll=412 and cc>=234 and cc<237) then grbp<="111";
	end if;
	if (ll=412 and cc>=238 and cc<241) then grbp<="111";
	end if;
	if (cc=8 and ll=413) then grbp<="111";
	end if;
	if (ll=413 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (ll=413 and cc>=22 and cc<24) then grbp<="111";
	end if;
	if (ll=413 and cc>=25 and cc<27) then grbp<="111";
	end if;
	if (cc=134 and ll=413) then grbp<="111";
	end if;
	if (cc=136 and ll=413) then grbp<="111";
	end if;
	if (cc=138 and ll=413) then grbp<="111";
	end if;
	if (cc=140 and ll=413) then grbp<="111";
	end if;
	if (ll=413 and cc>=140 and cc<142) then grbp<="111";
	end if;
	if (cc=148 and ll=413) then grbp<="111";
	end if;
	if (cc=151 and ll=413) then grbp<="111";
	end if;
	if (cc=155 and ll=413) then grbp<="111";
	end if;
	if (ll=413 and cc>=155 and cc<157) then grbp<="111";
	end if;
	if (cc=161 and ll=413) then grbp<="111";
	end if;
	if (ll=413 and cc>=161 and cc<163) then grbp<="111";
	end if;
	if (ll=413 and cc>=164 and cc<186) then grbp<="111";
	end if;
	if (cc=239 and ll=413) then grbp<="111";
	end if;
	if (cc=8 and ll=414) then grbp<="111";
	end if;
	if (ll=414 and cc>=8 and cc<14) then grbp<="111";
	end if;
	if (cc=140 and ll=414) then grbp<="111";
	end if;
	if (cc=164 and ll=414) then grbp<="111";
	end if;
	if (ll=414 and cc>=164 and cc<186) then grbp<="111";
	end if;
	if (ll=415 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (ll=415 and cc>=23 and cc<26) then grbp<="111";
	end if;
	if (cc=164 and ll=415) then grbp<="111";
	end if;
	if (ll=415 and cc>=164 and cc<186) then grbp<="111";
	end if;
	if (ll=416 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=25 and ll=416) then grbp<="111";
	end if;
	if (ll=416 and cc>=25 and cc<28) then grbp<="111";
	end if;
	if (ll=416 and cc>=164 and cc<186) then grbp<="111";
	end if;
	if (ll=417 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=62 and ll=417) then grbp<="111";
	end if;
	if (cc=164 and ll=417) then grbp<="111";
	end if;
	if (ll=417 and cc>=164 and cc<187) then grbp<="111";
	end if;
	if (ll=418 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (ll=418 and cc>=164 and cc<187) then grbp<="111";
	end if;
	if (ll=419 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=164 and ll=419) then grbp<="111";
	end if;
	if (ll=419 and cc>=164 and cc<166) then grbp<="111";
	end if;
	if (ll=419 and cc>=167 and cc<187) then grbp<="111";
	end if;
	if (ll=420 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=162 and ll=420) then grbp<="111";
	end if;
	if (ll=420 and cc>=162 and cc<187) then grbp<="111";
	end if;
	if (ll=421 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (ll=421 and cc>=165 and cc<187) then grbp<="111";
	end if;
	if (ll=422 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=26 and ll=422) then grbp<="111";
	end if;
	if (cc=164 and ll=422) then grbp<="111";
	end if;
	if (ll=422 and cc>=164 and cc<187) then grbp<="111";
	end if;
	if (ll=423 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=24 and ll=423) then grbp<="111";
	end if;
	if (cc=26 and ll=423) then grbp<="111";
	end if;
	if (cc=52 and ll=423) then grbp<="111";
	end if;
	if (cc=164 and ll=423) then grbp<="111";
	end if;
	if (ll=423 and cc>=164 and cc<188) then grbp<="111";
	end if;
	if (cc=8 and ll=424) then grbp<="111";
	end if;
	if (ll=424 and cc>=8 and cc<15) then grbp<="111";
	end if;
	if (cc=26 and ll=424) then grbp<="111";
	end if;
	if (ll=424 and cc>=26 and cc<28) then grbp<="111";
	end if;
	if (cc=163 and ll=424) then grbp<="111";
	end if;
	if (ll=424 and cc>=163 and cc<188) then grbp<="111";
	end if;
end if;
-------------------------------mode="100"--------------------clk---------------------
	 
if mode="100" then
    	 
	 -----------------------hour point------------CC + 5; LL + 13------RED "010"
	if cc<132 and cc>118 and ll<173 and ll>147 then grbp<="011";
	end if;

	if cc<132 and cc>119 and ll<53 and ll>27 then grbp<="010";
	end if;

	if cc<160 and cc>151 and ll<65 and ll>47 then grbp<="010";
	end if;

	if cc<181 and cc>172 and ll<109 and ll>91 then grbp<="010";
	end if;

	if cc<192 and cc>178 and ll<173 and ll>147 then grbp<="010";
	end if;

	if cc<181 and cc>172 and ll<229 and ll>211 then grbp<="010";
	end if;

	if cc<160 and cc>151 and ll<273 and ll>255 then grbp<="010";
	end if;

	if cc<132 and cc>119 and ll<293 and ll>267 then grbp<="010";
	end if;

	if cc<100 and cc>91 and ll<273 and ll>255 then grbp<="010";
	end if;

	if cc<78 and cc>69 and ll<229 and ll>211 then grbp<="010";
	end if;

	if cc<72 and cc>59 and ll<173 and ll>147 then grbp<="010";
	end if;

	if cc<77 and cc>68 and ll<109 and ll>91 then grbp<="010";
	end if;

	if cc<99 and cc>90 and ll<65 and ll>47 then grbp<="010";
	end if;

if ((PT0 ="0000" and PT1 ="0000") or (PT0 ="0001" and PT1 ="0010") or (PT0 ="0010" and PT1 ="0100")) then
	if ((cc=124 and ll>=128 and ll<167) or (cc=125 and ll>=106 and ll<167) or (cc=126 and ll>=139 and ll<167)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0001") or (PT0 ="0001" and PT1 ="0011")) then
	if ((cc=123 and ll>=162 and ll<166) or (cc=124 and ll>=158 and ll<167) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=151 and ll<163) or (cc=127 and ll>=150 and ll<159) or (cc=128 and ll>=146 and ll<156) or (cc=129 and ll>=143 and ll<152) or (cc=130 and ll>=140 and ll<149) or (cc=131 and ll>=136 and ll<146) or (cc=132 and ll>=133 and ll<138) or (cc=133 and ll>=131 and ll<134) or (cc=134 and ll>=127 and ll<131) or (cc=135 and ll>=124 and ll<127) or (cc=136 and ll>=120 and ll<124) or (cc=137 and ll>=117 and ll<120) or (cc=138 and ll>=113 and ll<117)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0010") or (PT0 ="0001" and PT1 ="0100")) then
	if ((cc=122 and ll>=161 and ll<164) or (cc=123 and ll>=160 and ll<166) or (cc=124 and ll>=158 and ll<165) or (cc=125 and ll>=157 and ll<164) or (cc=126 and ll>=156 and ll<163) or (cc=127 and ll>=155 and ll<161) or (cc=128 and ll>=154 and ll<160) or (cc=129 and ll>=153 and ll<159) or (cc=130 and ll>=153 and ll<158) or (cc=131 and ll>=152 and ll<157) or (cc=132 and ll>=151 and ll<156) or (cc=133 and ll>=149 and ll<154) or (cc=134 and ll>=148 and ll<153) or (cc=135 and ll>=147 and ll<152) or (cc=136 and ll>=146 and ll<148) or (cc=137 and ll>=145 and ll<147) or (cc=138 and ll>=144 and ll<146) or (cc=139 and ll>=143 and ll<145) or (cc=140 and ll>=142 and ll<144) or (cc=141 and ll>=141 and ll<143) or (cc=142 and ll=140) or (cc=143 and ll=139) or (cc=144 and ll>=137 and ll<139) or (cc=145 and ll>=136 and ll<138) or (cc=146 and ll>=135 and ll<137) or (cc=147 and ll>=134 and ll<136) or (cc=148 and ll=133)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0011") or (PT0 ="0001" and PT1 ="0101")) then
	if ((cc=122 and ll>=158 and ll<163) or (cc=123 and ll>=158 and ll<163) or (cc=124 and ll>=158 and ll<163) or (cc=125 and ll>=158 and ll<163) or (cc=126 and ll>=158 and ll<163) or (cc=127 and ll>=158 and ll<163) or (cc=128 and ll>=158 and ll<163) or (cc=129 and ll>=158 and ll<163) or (cc=130 and ll>=158 and ll<163) or (cc=131 and ll>=159 and ll<163) or (cc=132 and ll>=159 and ll<163) or (cc=133 and ll>=159 and ll<163) or (cc=134 and ll>=159 and ll<163) or (cc=135 and ll>=159 and ll<163) or (cc=136 and ll>=159 and ll<163) or (cc=137 and ll>=159 and ll<161) or (cc=138 and ll>=159 and ll<161) or (cc=139 and ll>=159 and ll<161) or (cc=140 and ll>=159 and ll<161) or (cc=141 and ll>=159 and ll<161) or (cc=142 and ll=160) or (cc=143 and ll=160) or (cc=144 and ll=160) or (cc=145 and ll=160) or (cc=146 and ll=160) or (cc=147 and ll=160) or (cc=148 and ll=160) or (cc=149 and ll=160) or (cc=150 and ll=160) or (cc=151 and ll=160) or (cc=152 and ll=160)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0100") or (PT0 ="0001" and PT1 ="0110")) then
	if ((cc=122 and ll>=157 and ll<160) or (cc=123 and ll>=155 and ll<161) or (cc=124 and ll>=156 and ll<162) or (cc=125 and ll>=157 and ll<164) or (cc=126 and ll>=159 and ll<165) or (cc=127 and ll>=160 and ll<166) or (cc=128 and ll>=161 and ll<167) or (cc=129 and ll>=162 and ll<168) or (cc=130 and ll>=163 and ll<169) or (cc=131 and ll>=166 and ll<171) or (cc=132 and ll>=167 and ll<172) or (cc=133 and ll>=168 and ll<173) or (cc=134 and ll>=169 and ll<173) or (cc=135 and ll>=170 and ll<173) or (cc=136 and ll>=171 and ll<174) or (cc=137 and ll>=172 and ll<175) or (cc=138 and ll>=174 and ll<176) or (cc=139 and ll>=175 and ll<177) or (cc=140 and ll=177) or (cc=141 and ll>=178 and ll<180) or (cc=142 and ll>=179 and ll<181) or (cc=143 and ll>=180 and ll<182) or (cc=144 and ll>=181 and ll<183) or (cc=145 and ll>=182 and ll<184) or (cc=146 and ll=184) or (cc=147 and ll=185) or (cc=148 and ll>=186 and ll<188)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0101") or (PT0 ="0001" and PT1 ="0111")) then
	if ((cc=123 and ll>=155 and ll<159) or (cc=124 and ll>=154 and ll<163) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=158 and ll<170) or (cc=127 and ll>=162 and ll<173) or (cc=128 and ll>=165 and ll<177) or (cc=129 and ll>=171 and ll<180) or (cc=130 and ll>=174 and ll<179) or (cc=131 and ll>=178 and ll<183) or (cc=132 and ll>=181 and ll<186) or (cc=133 and ll>=185 and ll<190) or (cc=134 and ll>=189 and ll<193) or (cc=135 and ll>=193 and ll<196) or (cc=136 and ll>=196 and ll<200) or (cc=137 and ll>=200 and ll<203) or (cc=138 and ll>=203 and ll<207) or (cc=139 and ll=207)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0110") or (PT0 ="0001" and PT1 ="1000")) then
	if ((cc=124 and ll>=154 and ll<182) or (cc=125 and ll>=154 and ll<215) or (cc=126 and ll>=154 and ll<193)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="0111") or (PT0 ="0001" and PT1 ="1001")) then
	if ((cc=112 and ll>=204 and ll<208) or (cc=113 and ll>=201 and ll<204) or (cc=114 and ll>=197 and ll<201) or (cc=115 and ll>=194 and ll<197) or (cc=116 and ll>=190 and ll<194) or (cc=117 and ll>=187 and ll<191) or (cc=118 and ll>=183 and ll<188) or (cc=119 and ll>=175 and ll<185) or (cc=120 and ll>=172 and ll<181) or (cc=121 and ll>=169 and ll<178) or (cc=122 and ll>=165 and ll<175) or (cc=123 and ll>=162 and ll<171) or (cc=124 and ll>=158 and ll<170) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=154 and ll<163) or (cc=127 and ll>=155 and ll<159)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="1000") or (PT0 ="0010" and PT1 ="0000")) then
	if ((cc=102 and ll=187) or (cc=103 and ll>=185 and ll<187) or (cc=104 and ll>=184 and ll<186) or (cc=105 and ll>=183 and ll<185) or (cc=106 and ll>=182 and ll<184) or (cc=107 and ll=181) or (cc=108 and ll=180) or (cc=109 and ll>=178 and ll<180) or (cc=110 and ll>=177 and ll<179) or (cc=111 and ll>=176 and ll<178) or (cc=112 and ll>=175 and ll<177) or (cc=113 and ll>=174 and ll<176) or (cc=114 and ll>=173 and ll<175) or (cc=115 and ll>=169 and ll<174) or (cc=116 and ll>=168 and ll<173) or (cc=117 and ll>=167 and ll<172) or (cc=118 and ll>=165 and ll<170) or (cc=119 and ll>=164 and ll<169) or (cc=120 and ll>=163 and ll<168) or (cc=121 and ll>=162 and ll<168) or (cc=122 and ll>=161 and ll<167) or (cc=123 and ll>=160 and ll<166) or (cc=124 and ll>=158 and ll<165) or (cc=125 and ll>=157 and ll<164) or (cc=126 and ll>=156 and ll<163) or (cc=127 and ll>=155 and ll<161) or (cc=128 and ll>=157 and ll<160)) then grbp<="111";
	end if;

elsif ((PT0 ="0000" and PT1 ="1001") or (PT0 ="0010" and PT1 ="0001")) then
	if ((cc=98 and ll=160) or (cc=99 and ll=160) or (cc=100 and ll=160) or (cc=101 and ll=160) or (cc=102 and ll=160) or (cc=103 and ll=160) or (cc=104 and ll=160) or (cc=105 and ll=160) or (cc=106 and ll=160) or (cc=107 and ll=160) or (cc=108 and ll=160) or (cc=109 and ll>=160 and ll<162) or (cc=110 and ll>=160 and ll<162) or (cc=111 and ll>=160 and ll<162) or (cc=112 and ll>=160 and ll<162) or (cc=113 and ll>=160 and ll<162) or (cc=114 and ll>=158 and ll<162) or (cc=115 and ll>=158 and ll<162) or (cc=116 and ll>=158 and ll<162) or (cc=117 and ll>=158 and ll<162) or (cc=118 and ll>=158 and ll<162) or (cc=119 and ll>=158 and ll<162) or (cc=120 and ll>=158 and ll<163) or (cc=121 and ll>=158 and ll<163) or (cc=122 and ll>=158 and ll<163) or (cc=123 and ll>=158 and ll<163) or (cc=124 and ll>=158 and ll<163) or (cc=125 and ll>=158 and ll<163) or (cc=126 and ll>=158 and ll<163) or (cc=127 and ll>=158 and ll<163) or (cc=128 and ll>=158 and ll<163)) then grbp<="111";
	end if;

elsif ((PT0 ="0001" and PT1 ="0000") or (PT0 ="0010" and PT1 ="0010")) then
	if ((cc=102 and ll>=133 and ll<135) or (cc=103 and ll=135) or (cc=104 and ll=136) or (cc=105 and ll>=137 and ll<139) or (cc=106 and ll>=138 and ll<140) or (cc=107 and ll>=139 and ll<141) or (cc=108 and ll>=140 and ll<142) or (cc=109 and ll>=141 and ll<143) or (cc=110 and ll=143) or (cc=111 and ll>=144 and ll<146) or (cc=112 and ll>=145 and ll<147) or (cc=113 and ll>=146 and ll<149) or (cc=114 and ll>=147 and ll<150) or (cc=115 and ll>=148 and ll<151) or (cc=116 and ll>=148 and ll<152) or (cc=117 and ll>=148 and ll<153) or (cc=118 and ll>=149 and ll<154) or (cc=119 and ll>=150 and ll<155) or (cc=120 and ll>=152 and ll<158) or (cc=121 and ll>=153 and ll<159) or (cc=122 and ll>=154 and ll<160) or (cc=123 and ll>=155 and ll<161) or (cc=124 and ll>=156 and ll<162) or (cc=125 and ll>=157 and ll<164) or (cc=126 and ll>=159 and ll<165) or (cc=127 and ll>=160 and ll<166) or (cc=128 and ll>=161 and ll<164)) then grbp<="111";
	end if;

elsif ((PT0 ="0001" and PT1 ="0001") or (PT0 ="0010" and PT1 ="0011")) then
	if ((cc=111 and ll=113) or (cc=112 and ll>=114 and ll<118) or (cc=113 and ll>=118 and ll<121) or (cc=114 and ll>=121 and ll<125) or (cc=115 and ll>=125 and ll<128) or (cc=116 and ll>=128 and ll<132) or (cc=117 and ll>=131 and ll<136) or (cc=118 and ll>=135 and ll<140) or (cc=119 and ll>=138 and ll<143) or (cc=120 and ll>=142 and ll<147) or (cc=121 and ll>=141 and ll<150) or (cc=122 and ll>=144 and ll<156) or (cc=123 and ll>=148 and ll<159) or (cc=124 and ll>=151 and ll<163) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=158 and ll<167) or (cc=127 and ll>=162 and ll<166)) then grbp<="111";
	end if;


end if;
	if cc<134 and cc>129 and ll<46 and ll>36 then grbp<="010";
	end if;

	if cc<140 and cc>135 and ll<48 and ll>38 then grbp<="010";
	end if;

	if cc<146 and cc>141 and ll<51 and ll>41 then grbp<="010";
	end if;

	if cc<152 and cc>147 and ll<55 and ll>45 then grbp<="010";
	end if;

	if cc<163 and cc>158 and ll<68 and ll>58 then grbp<="010";
	end if;

	if cc<168 and cc>163 and ll<76 and ll>66 then grbp<="010";
	end if;

	if cc<172 and cc>167 and ll<85 and ll>75 then grbp<="010";
	end if;

	if cc<176 and cc>171 and ll<94 and ll>84 then grbp<="010";
	end if;

	if cc<182 and cc>177 and ll<116 and ll>106 then grbp<="010";
	end if;

	if cc<185 and cc>180 and ll<128 and ll>118 then grbp<="010";
	end if;

	if cc<186 and cc>181 and ll<140 and ll>130 then grbp<="010";
	end if;

	if cc<187 and cc>182 and ll<152 and ll>142 then grbp<="010";
	end if;

	if cc<187 and cc>182 and ll<178 and ll>168 then grbp<="010";
	end if;

	if cc<186 and cc>181 and ll<190 and ll>180 then grbp<="010";
	end if;

	if cc<185 and cc>180 and ll<202 and ll>192 then grbp<="010";
	end if;

	if cc<182 and cc>177 and ll<214 and ll>204 then grbp<="010";
	end if;

	if cc<176 and cc>171 and ll<236 and ll>226 then grbp<="010";
	end if;

	if cc<172 and cc>167 and ll<245 and ll>235 then grbp<="010";
	end if;

	if cc<168 and cc>163 and ll<254 and ll>244 then grbp<="010";
	end if;

	if cc<163 and cc>158 and ll<262 and ll>252 then grbp<="010";
	end if;

	if cc<152 and cc>147 and ll<275 and ll>265 then grbp<="010";
	end if;

	if cc<146 and cc>141 and ll<279 and ll>269 then grbp<="010";
	end if;

	if cc<140 and cc>135 and ll<282 and ll>272 then grbp<="010";
	end if;

	if cc<134 and cc>129 and ll<284 and ll>274 then grbp<="010";
	end if;

	if cc<121 and cc>116 and ll<284 and ll>274 then grbp<="010";
	end if;

	if cc<115 and cc>110 and ll<282 and ll>272 then grbp<="010";
	end if;

	if cc<109 and cc>104 and ll<279 and ll>269 then grbp<="010";
	end if;

	if cc<103 and cc>98 and ll<275 and ll>265 then grbp<="010";
	end if;

	if cc<92 and cc>87 and ll<262 and ll>252 then grbp<="010";
	end if;

	if cc<87 and cc>82 and ll<254 and ll>244 then grbp<="010";
	end if;

	if cc<83 and cc>78 and ll<245 and ll>235 then grbp<="010";
	end if;

	if cc<79 and cc>74 and ll<236 and ll>226 then grbp<="010";
	end if;

	if cc<73 and cc>68 and ll<214 and ll>204 then grbp<="010";
	end if;

	if cc<70 and cc>65 and ll<202 and ll>192 then grbp<="010";
	end if;

	if cc<69 and cc>64 and ll<190 and ll>180 then grbp<="010";
	end if;

	if cc<68 and cc>63 and ll<178 and ll>168 then grbp<="010";
	end if;

	if cc<68 and cc>63 and ll<153 and ll>143 then grbp<="010";
	end if;

	if cc<69 and cc>64 and ll<140 and ll>130 then grbp<="010";
	end if;

	if cc<70 and cc>65 and ll<128 and ll>118 then grbp<="010";
	end if;

	if cc<73 and cc>68 and ll<116 and ll>106 then grbp<="010";
	end if;

	if cc<79 and cc>74 and ll<95 and ll>85 then grbp<="010";
	end if;

	if cc<83 and cc>78 and ll<85 and ll>75 then grbp<="010";
	end if;

	if cc<87 and cc>82 and ll<76 and ll>66 then grbp<="010";
	end if;

	if cc<92 and cc>87 and ll<68 and ll>58 then grbp<="010";
	end if;

	if cc<103 and cc>98 and ll<55 and ll>45 then grbp<="010";
	end if;

	if cc<109 and cc>104 and ll<51 and ll>41 then grbp<="010";
	end if;

	if cc<115 and cc>110 and ll<48 and ll>38 then grbp<="010";
	end if;

	if cc<121 and cc>116 and ll<46 and ll>36 then grbp<="010";
	end if;

if ((PT2 ="0000" and PT3 ="0000")) then
	if ((cc=123 and ll>=146 and ll<160) or (cc=124 and ll>=102 and ll<169) or (cc=125 and ll>=80 and ll<169) or (cc=126 and ll>=113 and ll<169) or (cc=127 and ll>=157 and ll<169)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0001")) then
	if ((cc=123 and ll>=161 and ll<169) or (cc=124 and ll>=146 and ll<169) or (cc=125 and ll>=131 and ll<169) or (cc=126 and ll>=122 and ll<169) or (cc=127 and ll>=102 and ll<169) or (cc=128 and ll>=92 and ll<131) or (cc=129 and ll>=80 and ll<92)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0010")) then
	if ((cc=123 and ll>=160 and ll<168) or (cc=124 and ll>=151 and ll<169) or (cc=125 and ll>=146 and ll<169) or (cc=126 and ll>=136 and ll<170) or (cc=127 and ll>=127 and ll<166) or (cc=128 and ll>=123 and ll<147) or (cc=129 and ll>=113 and ll<137) or (cc=130 and ll>=103 and ll<127) or (cc=131 and ll>=98 and ll<118) or (cc=132 and ll>=90 and ll<98) or (cc=133 and ll>=82 and ll<90)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0011")) then
	if ((cc=122 and ll>=166 and ll<168) or (cc=123 and ll>=160 and ll<168) or (cc=124 and ll>=153 and ll<169) or (cc=125 and ll>=148 and ll<169) or (cc=126 and ll>=145 and ll<170) or (cc=127 and ll>=138 and ll<164) or (cc=128 and ll>=133 and ll<151) or (cc=129 and ll>=126 and ll<145) or (cc=130 and ll>=124 and ll<139) or (cc=131 and ll>=117 and ll<133) or (cc=132 and ll>=111 and ll<126) or (cc=133 and ll>=105 and ll<121) or (cc=134 and ll>=102 and ll<108) or (cc=135 and ll>=95 and ll<102) or (cc=136 and ll>=90 and ll<95) or (cc=137 and ll>=84 and ll<90)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0100")) then
	if ((cc=122 and ll>=164 and ll<168) or (cc=123 and ll>=160 and ll<168) or (cc=124 and ll>=155 and ll<169) or (cc=125 and ll>=151 and ll<170) or (cc=126 and ll>=146 and ll<168) or (cc=127 and ll>=145 and ll<164) or (cc=128 and ll>=140 and ll<154) or (cc=129 and ll>=135 and ll<150) or (cc=130 and ll>=131 and ll<145) or (cc=131 and ll>=126 and ll<141) or (cc=132 and ll>=124 and ll<136) or (cc=133 and ll>=119 and ll<132) or (cc=134 and ll>=115 and ll<127) or (cc=135 and ll>=110 and ll<122) or (cc=136 and ll>=107 and ll<113) or (cc=137 and ll>=104 and ll<109) or (cc=138 and ll>=100 and ll<104) or (cc=139 and ll>=95 and ll<100) or (cc=140 and ll>=91 and ll<95) or (cc=141 and ll>=87 and ll<91)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0101")) then
	if ((cc=122 and ll>=163 and ll<167) or (cc=123 and ll>=159 and ll<168) or (cc=124 and ll>=156 and ll<169) or (cc=125 and ll>=152 and ll<170) or (cc=126 and ll>=149 and ll<166) or (cc=127 and ll>=146 and ll<163) or (cc=128 and ll>=144 and ll<156) or (cc=129 and ll>=141 and ll<152) or (cc=130 and ll>=137 and ll<149) or (cc=131 and ll>=134 and ll<146) or (cc=132 and ll>=130 and ll<142) or (cc=133 and ll>=128 and ll<139) or (cc=134 and ll>=126 and ll<135) or (cc=135 and ll>=122 and ll<132) or (cc=136 and ll>=119 and ll<128) or (cc=137 and ll>=115 and ll<125) or (cc=138 and ll>=112 and ll<121) or (cc=139 and ll>=109 and ll<113) or (cc=140 and ll>=106 and ll<110) or (cc=141 and ll>=103 and ll<106) or (cc=142 and ll>=99 and ll<103) or (cc=143 and ll>=96 and ll<99) or (cc=144 and ll>=92 and ll<96) or (cc=145 and ll>=91 and ll<93)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0110")) then
	if ((cc=121 and ll=165) or (cc=122 and ll>=162 and ll<167) or (cc=123 and ll>=159 and ll<169) or (cc=124 and ll>=157 and ll<170) or (cc=125 and ll>=154 and ll<169) or (cc=126 and ll>=151 and ll<166) or (cc=127 and ll>=149 and ll<163) or (cc=128 and ll>=147 and ll<157) or (cc=129 and ll>=144 and ll<154) or (cc=130 and ll>=142 and ll<152) or (cc=131 and ll>=139 and ll<149) or (cc=132 and ll>=136 and ll<146) or (cc=133 and ll>=134 and ll<144) or (cc=134 and ll>=130 and ll<140) or (cc=135 and ll>=129 and ll<138) or (cc=136 and ll>=127 and ll<135) or (cc=137 and ll>=124 and ll<132) or (cc=138 and ll>=121 and ll<130) or (cc=139 and ll>=119 and ll<127) or (cc=140 and ll>=116 and ll<124) or (cc=141 and ll>=113 and ll<118) or (cc=142 and ll>=112 and ll<115) or (cc=143 and ll>=109 and ll<112) or (cc=144 and ll>=107 and ll<109) or (cc=145 and ll>=104 and ll<107) or (cc=146 and ll>=101 and ll<104) or (cc=147 and ll>=98 and ll<101) or (cc=148 and ll>=95 and ll<99)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="0111")) then
	if ((cc=121 and ll=164) or (cc=122 and ll>=162 and ll<167) or (cc=123 and ll>=159 and ll<168) or (cc=124 and ll>=157 and ll<170) or (cc=125 and ll>=155 and ll<167) or (cc=126 and ll>=153 and ll<165) or (cc=127 and ll>=151 and ll<163) or (cc=128 and ll>=148 and ll<158) or (cc=129 and ll>=147 and ll<156) or (cc=130 and ll>=145 and ll<153) or (cc=131 and ll>=143 and ll<151) or (cc=132 and ll>=141 and ll<149) or (cc=133 and ll>=139 and ll<147) or (cc=134 and ll>=136 and ll<144) or (cc=135 and ll>=134 and ll<142) or (cc=136 and ll>=132 and ll<140) or (cc=137 and ll>=131 and ll<138) or (cc=138 and ll>=129 and ll<136) or (cc=139 and ll>=127 and ll<133) or (cc=140 and ll>=124 and ll<131) or (cc=141 and ll>=122 and ll<129) or (cc=142 and ll>=120 and ll<124) or (cc=143 and ll>=118 and ll<122) or (cc=144 and ll>=116 and ll<119) or (cc=145 and ll>=115 and ll<117) or (cc=146 and ll>=112 and ll<115) or (cc=147 and ll>=110 and ll<113) or (cc=148 and ll>=108 and ll<110) or (cc=149 and ll>=106 and ll<108) or (cc=150 and ll>=103 and ll<106) or (cc=151 and ll>=101 and ll<104) or (cc=152 and ll=100)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="1000")) then
	if ((cc=121 and ll>=162 and ll<165) or (cc=122 and ll>=161 and ll<166) or (cc=123 and ll>=159 and ll<169) or (cc=124 and ll>=157 and ll<169) or (cc=125 and ll>=155 and ll<167) or (cc=126 and ll>=154 and ll<165) or (cc=127 and ll>=152 and ll<163) or (cc=128 and ll>=150 and ll<159) or (cc=129 and ll>=148 and ll<157) or (cc=130 and ll>=148 and ll<155) or (cc=131 and ll>=146 and ll<153) or (cc=132 and ll>=144 and ll<152) or (cc=133 and ll>=142 and ll<150) or (cc=134 and ll>=140 and ll<148) or (cc=135 and ll>=138 and ll<146) or (cc=136 and ll>=137 and ll<144) or (cc=137 and ll>=135 and ll<142) or (cc=138 and ll>=134 and ll<141) or (cc=139 and ll>=133 and ll<139) or (cc=140 and ll>=131 and ll<137) or (cc=141 and ll>=129 and ll<136) or (cc=142 and ll>=127 and ll<134) or (cc=143 and ll>=126 and ll<132) or (cc=144 and ll>=124 and ll<127) or (cc=145 and ll>=122 and ll<125) or (cc=146 and ll>=120 and ll<123) or (cc=147 and ll>=120 and ll<122) or (cc=148 and ll>=118 and ll<120) or (cc=149 and ll>=116 and ll<118) or (cc=150 and ll>=114 and ll<116) or (cc=151 and ll>=112 and ll<115) or (cc=152 and ll>=110 and ll<113) or (cc=153 and ll>=109 and ll<111) or (cc=154 and ll>=107 and ll<109) or (cc=155 and ll=106)) then grbp<="001";
	end if;

elsif ((PT2 ="0000" and PT3 ="1001")) then
	if ((cc=121 and ll>=162 and ll<165) or (cc=122 and ll>=161 and ll<167) or (cc=123 and ll>=159 and ll<169) or (cc=124 and ll>=158 and ll<168) or (cc=125 and ll>=156 and ll<167) or (cc=126 and ll>=155 and ll<165) or (cc=127 and ll>=153 and ll<164) or (cc=128 and ll>=152 and ll<160) or (cc=129 and ll>=150 and ll<158) or (cc=130 and ll>=149 and ll<157) or (cc=131 and ll>=148 and ll<155) or (cc=132 and ll>=147 and ll<154) or (cc=133 and ll>=145 and ll<152) or (cc=134 and ll>=144 and ll<151) or (cc=135 and ll>=142 and ll<149) or (cc=136 and ll>=141 and ll<148) or (cc=137 and ll>=140 and ll<146) or (cc=138 and ll>=138 and ll<145) or (cc=139 and ll>=137 and ll<144) or (cc=140 and ll>=136 and ll<142) or (cc=141 and ll>=135 and ll<141) or (cc=142 and ll>=133 and ll<139) or (cc=143 and ll>=132 and ll<138) or (cc=144 and ll>=130 and ll<136) or (cc=145 and ll>=129 and ll<135) or (cc=146 and ll>=128 and ll<131) or (cc=147 and ll>=126 and ll<129) or (cc=148 and ll>=125 and ll<128) or (cc=149 and ll=125) or (cc=150 and ll>=123 and ll<125) or (cc=151 and ll=122) or (cc=152 and ll>=120 and ll<122) or (cc=153 and ll=119) or (cc=154 and ll>=117 and ll<119) or (cc=155 and ll=116) or (cc=156 and ll=115) or (cc=157 and ll>=113 and ll<115)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0000")) then
	if ((cc=121 and ll>=161 and ll<164) or (cc=122 and ll>=160 and ll<167) or (cc=123 and ll>=158 and ll<168) or (cc=124 and ll>=157 and ll<167) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=155 and ll<165) or (cc=127 and ll>=154 and ll<163) or (cc=128 and ll>=153 and ll<160) or (cc=129 and ll>=151 and ll<159) or (cc=130 and ll>=150 and ll<158) or (cc=131 and ll>=150 and ll<157) or (cc=132 and ll>=149 and ll<156) or (cc=133 and ll>=148 and ll<154) or (cc=134 and ll>=147 and ll<153) or (cc=135 and ll>=146 and ll<152) or (cc=136 and ll>=145 and ll<151) or (cc=137 and ll>=143 and ll<150) or (cc=138 and ll>=142 and ll<149) or (cc=139 and ll>=141 and ll<147) or (cc=140 and ll>=140 and ll<146) or (cc=141 and ll>=140 and ll<145) or (cc=142 and ll>=139 and ll<144) or (cc=143 and ll>=138 and ll<143) or (cc=144 and ll>=137 and ll<142) or (cc=145 and ll>=136 and ll<141) or (cc=146 and ll>=134 and ll<139) or (cc=147 and ll>=133 and ll<136) or (cc=148 and ll>=132 and ll<134) or (cc=149 and ll>=131 and ll<133) or (cc=150 and ll>=130 and ll<132) or (cc=151 and ll>=129 and ll<131) or (cc=152 and ll>=128 and ll<130) or (cc=153 and ll>=127 and ll<129) or (cc=154 and ll>=126 and ll<128) or (cc=155 and ll=125) or (cc=156 and ll=124) or (cc=157 and ll>=122 and ll<124) or (cc=158 and ll>=121 and ll<123) or (cc=159 and ll>=120 and ll<122) or (cc=160 and ll=120)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0001")) then
	if ((cc=121 and ll>=160 and ll<164) or (cc=122 and ll>=159 and ll<168) or (cc=123 and ll>=158 and ll<168) or (cc=124 and ll>=157 and ll<167) or (cc=125 and ll>=156 and ll<165) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=155 and ll<164) or (cc=128 and ll>=154 and ll<161) or (cc=129 and ll>=153 and ll<160) or (cc=130 and ll>=152 and ll<159) or (cc=131 and ll>=152 and ll<158) or (cc=132 and ll>=151 and ll<157) or (cc=133 and ll>=150 and ll<156) or (cc=134 and ll>=150 and ll<155) or (cc=135 and ll>=149 and ll<155) or (cc=136 and ll>=148 and ll<153) or (cc=137 and ll>=147 and ll<153) or (cc=138 and ll>=146 and ll<152) or (cc=139 and ll>=145 and ll<151) or (cc=140 and ll>=144 and ll<150) or (cc=141 and ll>=143 and ll<149) or (cc=142 and ll>=144 and ll<148) or (cc=143 and ll>=143 and ll<147) or (cc=144 and ll>=142 and ll<146) or (cc=145 and ll>=141 and ll<146) or (cc=146 and ll>=140 and ll<144) or (cc=147 and ll>=139 and ll<144) or (cc=148 and ll>=138 and ll<141) or (cc=149 and ll>=137 and ll<140) or (cc=150 and ll>=136 and ll<139) or (cc=151 and ll>=135 and ll<138) or (cc=152 and ll>=135 and ll<137) or (cc=153 and ll=135) or (cc=154 and ll=134) or (cc=155 and ll=133) or (cc=156 and ll>=132 and ll<134) or (cc=157 and ll=131) or (cc=158 and ll>=130 and ll<132) or (cc=159 and ll>=129 and ll<131) or (cc=160 and ll=129) or (cc=161 and ll=128) or (cc=162 and ll=127)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0010")) then
	if ((cc=121 and ll>=159 and ll<163) or (cc=122 and ll>=159 and ll<167) or (cc=123 and ll>=158 and ll<167) or (cc=124 and ll>=157 and ll<166) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=155 and ll<164) or (cc=128 and ll>=155 and ll<161) or (cc=129 and ll>=154 and ll<161) or (cc=130 and ll>=153 and ll<160) or (cc=131 and ll>=153 and ll<159) or (cc=132 and ll>=153 and ll<159) or (cc=133 and ll>=152 and ll<158) or (cc=134 and ll>=152 and ll<157) or (cc=135 and ll>=151 and ll<157) or (cc=136 and ll>=151 and ll<156) or (cc=137 and ll>=150 and ll<155) or (cc=138 and ll>=149 and ll<155) or (cc=139 and ll>=148 and ll<154) or (cc=140 and ll>=148 and ll<154) or (cc=141 and ll>=147 and ll<153) or (cc=142 and ll>=147 and ll<152) or (cc=143 and ll>=147 and ll<151) or (cc=144 and ll>=146 and ll<151) or (cc=145 and ll>=146 and ll<150) or (cc=146 and ll>=145 and ll<150) or (cc=147 and ll>=144 and ll<149) or (cc=148 and ll>=144 and ll<148) or (cc=149 and ll>=143 and ll<145) or (cc=150 and ll>=143 and ll<145) or (cc=151 and ll>=142 and ll<144) or (cc=152 and ll>=141 and ll<144) or (cc=153 and ll=142) or (cc=154 and ll=141) or (cc=155 and ll=140) or (cc=156 and ll>=139 and ll<141) or (cc=157 and ll=139) or (cc=158 and ll>=138 and ll<140) or (cc=159 and ll=138) or (cc=160 and ll=137) or (cc=161 and ll>=136 and ll<138) or (cc=162 and ll=136) or (cc=163 and ll=135)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0011")) then
	if ((cc=121 and ll>=159 and ll<165) or (cc=122 and ll>=158 and ll<167) or (cc=123 and ll>=158 and ll<166) or (cc=124 and ll>=157 and ll<166) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=156 and ll<164) or (cc=128 and ll>=156 and ll<162) or (cc=129 and ll>=155 and ll<161) or (cc=130 and ll>=155 and ll<161) or (cc=131 and ll>=154 and ll<161) or (cc=132 and ll>=154 and ll<160) or (cc=133 and ll>=154 and ll<160) or (cc=134 and ll>=154 and ll<159) or (cc=135 and ll>=154 and ll<159) or (cc=136 and ll>=153 and ll<158) or (cc=137 and ll>=153 and ll<158) or (cc=138 and ll>=152 and ll<157) or (cc=139 and ll>=152 and ll<157) or (cc=140 and ll>=151 and ll<157) or (cc=141 and ll>=151 and ll<156) or (cc=142 and ll>=150 and ll<156) or (cc=143 and ll>=151 and ll<155) or (cc=144 and ll>=151 and ll<155) or (cc=145 and ll>=150 and ll<155) or (cc=146 and ll>=150 and ll<154) or (cc=147 and ll>=149 and ll<154) or (cc=148 and ll>=149 and ll<153) or (cc=149 and ll>=149 and ll<151) or (cc=150 and ll>=148 and ll<150) or (cc=151 and ll>=148 and ll<150) or (cc=152 and ll>=147 and ll<149) or (cc=153 and ll>=147 and ll<149) or (cc=154 and ll>=147 and ll<149) or (cc=155 and ll=147) or (cc=156 and ll=147) or (cc=157 and ll=146) or (cc=158 and ll=146) or (cc=159 and ll>=145 and ll<147) or (cc=160 and ll=145) or (cc=161 and ll>=144 and ll<146) or (cc=162 and ll=144) or (cc=163 and ll=144) or (cc=164 and ll=143)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0100")) then
	if ((cc=121 and ll>=158 and ll<166) or (cc=122 and ll>=158 and ll<166) or (cc=123 and ll>=157 and ll<166) or (cc=124 and ll>=157 and ll<165) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=157 and ll<165) or (cc=127 and ll>=156 and ll<165) or (cc=128 and ll>=156 and ll<162) or (cc=129 and ll>=156 and ll<162) or (cc=130 and ll>=156 and ll<162) or (cc=131 and ll>=156 and ll<162) or (cc=132 and ll>=156 and ll<162) or (cc=133 and ll>=156 and ll<161) or (cc=134 and ll>=156 and ll<161) or (cc=135 and ll>=156 and ll<161) or (cc=136 and ll>=156 and ll<161) or (cc=137 and ll>=155 and ll<161) or (cc=138 and ll>=155 and ll<160) or (cc=139 and ll>=155 and ll<160) or (cc=140 and ll>=155 and ll<160) or (cc=141 and ll>=154 and ll<160) or (cc=142 and ll>=154 and ll<159) or (cc=143 and ll>=154 and ll<159) or (cc=144 and ll>=155 and ll<159) or (cc=145 and ll>=155 and ll<159) or (cc=146 and ll>=154 and ll<159) or (cc=147 and ll>=154 and ll<158) or (cc=148 and ll>=154 and ll<158) or (cc=149 and ll>=154 and ll<156) or (cc=150 and ll>=154 and ll<156) or (cc=151 and ll>=153 and ll<155) or (cc=152 and ll>=153 and ll<155) or (cc=153 and ll>=153 and ll<155) or (cc=154 and ll>=153 and ll<155) or (cc=155 and ll>=153 and ll<155) or (cc=156 and ll=153) or (cc=157 and ll=153) or (cc=158 and ll=153) or (cc=159 and ll=153) or (cc=160 and ll>=152 and ll<154) or (cc=161 and ll=152) or (cc=162 and ll=152) or (cc=163 and ll=152) or (cc=164 and ll=152) or (cc=165 and ll=151)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0101")) then
	if ((cc=121 and ll>=157 and ll<165) or (cc=122 and ll>=157 and ll<165) or (cc=123 and ll>=157 and ll<165) or (cc=124 and ll>=157 and ll<165) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=157 and ll<165) or (cc=127 and ll>=157 and ll<165) or (cc=128 and ll>=157 and ll<163) or (cc=129 and ll>=157 and ll<163) or (cc=130 and ll>=157 and ll<163) or (cc=131 and ll>=157 and ll<163) or (cc=132 and ll>=157 and ll<163) or (cc=133 and ll>=158 and ll<163) or (cc=134 and ll>=158 and ll<163) or (cc=135 and ll>=158 and ll<163) or (cc=136 and ll>=158 and ll<163) or (cc=137 and ll>=158 and ll<163) or (cc=138 and ll>=158 and ll<163) or (cc=139 and ll>=158 and ll<163) or (cc=140 and ll>=158 and ll<163) or (cc=141 and ll>=158 and ll<163) or (cc=142 and ll>=158 and ll<163) or (cc=143 and ll>=158 and ll<163) or (cc=144 and ll>=159 and ll<163) or (cc=145 and ll>=159 and ll<163) or (cc=146 and ll>=159 and ll<163) or (cc=147 and ll>=159 and ll<163) or (cc=148 and ll>=159 and ll<163) or (cc=149 and ll>=159 and ll<163) or (cc=150 and ll>=159 and ll<161) or (cc=151 and ll>=159 and ll<161) or (cc=152 and ll>=159 and ll<161) or (cc=153 and ll>=159 and ll<161) or (cc=154 and ll>=159 and ll<161) or (cc=155 and ll=160) or (cc=156 and ll=160) or (cc=157 and ll=160) or (cc=158 and ll=160) or (cc=159 and ll=160) or (cc=160 and ll=160) or (cc=161 and ll=160) or (cc=162 and ll=160) or (cc=163 and ll=160) or (cc=164 and ll=160) or (cc=165 and ll=160)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0110")) then
	if ((cc=121 and ll>=156 and ll<164) or (cc=122 and ll>=156 and ll<164) or (cc=123 and ll>=157 and ll<165) or (cc=124 and ll>=157 and ll<165) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=157 and ll<165) or (cc=127 and ll>=157 and ll<164) or (cc=128 and ll>=158 and ll<164) or (cc=129 and ll>=158 and ll<164) or (cc=130 and ll>=158 and ll<164) or (cc=131 and ll>=158 and ll<164) or (cc=132 and ll>=158 and ll<165) or (cc=133 and ll>=160 and ll<165) or (cc=134 and ll>=160 and ll<165) or (cc=135 and ll>=160 and ll<165) or (cc=136 and ll>=160 and ll<165) or (cc=137 and ll>=160 and ll<166) or (cc=138 and ll>=161 and ll<166) or (cc=139 and ll>=161 and ll<166) or (cc=140 and ll>=161 and ll<166) or (cc=141 and ll>=161 and ll<166) or (cc=142 and ll>=161 and ll<167) or (cc=143 and ll>=162 and ll<167) or (cc=144 and ll>=163 and ll<167) or (cc=145 and ll>=163 and ll<167) or (cc=146 and ll>=163 and ll<167) or (cc=147 and ll>=163 and ll<168) or (cc=148 and ll>=164 and ll<168) or (cc=149 and ll>=164 and ll<166) or (cc=150 and ll>=164 and ll<166) or (cc=151 and ll>=164 and ll<166) or (cc=152 and ll>=165 and ll<167) or (cc=153 and ll>=165 and ll<167) or (cc=154 and ll>=165 and ll<167) or (cc=155 and ll=166) or (cc=156 and ll=166) or (cc=157 and ll=167) or (cc=158 and ll=167) or (cc=159 and ll=167) or (cc=160 and ll=167) or (cc=161 and ll=167) or (cc=162 and ll=168) or (cc=163 and ll=168) or (cc=164 and ll=168) or (cc=165 and ll=168)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="0111")) then
	if ((cc=121 and ll>=155 and ll<163) or (cc=122 and ll>=156 and ll<164) or (cc=123 and ll>=156 and ll<164) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=157 and ll<166) or (cc=127 and ll>=158 and ll<164) or (cc=128 and ll>=158 and ll<164) or (cc=129 and ll>=159 and ll<165) or (cc=130 and ll>=159 and ll<165) or (cc=131 and ll>=159 and ll<166) or (cc=132 and ll>=160 and ll<166) or (cc=133 and ll>=161 and ll<166) or (cc=134 and ll>=162 and ll<167) or (cc=135 and ll>=162 and ll<167) or (cc=136 and ll>=163 and ll<168) or (cc=137 and ll>=163 and ll<168) or (cc=138 and ll>=163 and ll<169) or (cc=139 and ll>=164 and ll<169) or (cc=140 and ll>=164 and ll<170) or (cc=141 and ll>=165 and ll<170) or (cc=142 and ll>=165 and ll<170) or (cc=143 and ll>=165 and ll<171) or (cc=144 and ll>=167 and ll<171) or (cc=145 and ll>=167 and ll<172) or (cc=146 and ll>=168 and ll<172) or (cc=147 and ll>=168 and ll<172) or (cc=148 and ll>=168 and ll<173) or (cc=149 and ll>=169 and ll<171) or (cc=150 and ll>=169 and ll<172) or (cc=151 and ll>=170 and ll<172) or (cc=152 and ll>=170 and ll<173) or (cc=153 and ll>=171 and ll<173) or (cc=154 and ll=172) or (cc=155 and ll=173) or (cc=156 and ll=173) or (cc=157 and ll>=173 and ll<175) or (cc=158 and ll=174) or (cc=159 and ll=174) or (cc=160 and ll=175) or (cc=161 and ll=175) or (cc=162 and ll>=175 and ll<177) or (cc=163 and ll=176) or (cc=164 and ll=176)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="1000")) then
	if ((cc=121 and ll>=156 and ll<163) or (cc=122 and ll>=155 and ll<164) or (cc=123 and ll>=155 and ll<164) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=157 and ll<165) or (cc=126 and ll>=157 and ll<166) or (cc=127 and ll>=158 and ll<164) or (cc=128 and ll>=159 and ll<165) or (cc=129 and ll>=159 and ll<166) or (cc=130 and ll>=160 and ll<167) or (cc=131 and ll>=161 and ll<167) or (cc=132 and ll>=161 and ll<168) or (cc=133 and ll>=163 and ll<168) or (cc=134 and ll>=164 and ll<169) or (cc=135 and ll>=164 and ll<170) or (cc=136 and ll>=165 and ll<170) or (cc=137 and ll>=165 and ll<171) or (cc=138 and ll>=166 and ll<172) or (cc=139 and ll>=167 and ll<172) or (cc=140 and ll>=167 and ll<173) or (cc=141 and ll>=168 and ll<174) or (cc=142 and ll>=169 and ll<174) or (cc=143 and ll>=170 and ll<175) or (cc=144 and ll>=171 and ll<175) or (cc=145 and ll>=172 and ll<176) or (cc=146 and ll>=172 and ll<177) or (cc=147 and ll>=173 and ll<177) or (cc=148 and ll>=173 and ll<176) or (cc=149 and ll>=174 and ll<177) or (cc=150 and ll>=175 and ll<177) or (cc=151 and ll>=176 and ll<178) or (cc=152 and ll>=176 and ll<178) or (cc=153 and ll>=177 and ll<179) or (cc=154 and ll>=178 and ll<180) or (cc=155 and ll>=179 and ll<181) or (cc=156 and ll=180) or (cc=157 and ll=181) or (cc=158 and ll=181) or (cc=159 and ll=182) or (cc=160 and ll>=182 and ll<184) or (cc=161 and ll=183) or (cc=162 and ll=184) or (cc=163 and ll>=184 and ll<186)) then grbp<="001";
	end if;

elsif ((PT2 ="0001" and PT3 ="1001")) then
	if ((cc=121 and ll>=157 and ll<162) or (cc=122 and ll>=154 and ll<163) or (cc=123 and ll>=155 and ll<164) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=156 and ll<165) or (cc=126 and ll>=157 and ll<166) or (cc=127 and ll>=158 and ll<165) or (cc=128 and ll>=159 and ll<166) or (cc=129 and ll>=160 and ll<167) or (cc=130 and ll>=161 and ll<168) or (cc=131 and ll>=162 and ll<169) or (cc=132 and ll>=163 and ll<170) or (cc=133 and ll>=165 and ll<171) or (cc=134 and ll>=165 and ll<171) or (cc=135 and ll>=166 and ll<172) or (cc=136 and ll>=167 and ll<173) or (cc=137 and ll>=168 and ll<174) or (cc=138 and ll>=169 and ll<175) or (cc=139 and ll>=170 and ll<176) or (cc=140 and ll>=171 and ll<177) or (cc=141 and ll>=172 and ll<177) or (cc=142 and ll>=173 and ll<179) or (cc=143 and ll>=174 and ll<179) or (cc=144 and ll>=176 and ll<180) or (cc=145 and ll>=176 and ll<181) or (cc=146 and ll>=177 and ll<182) or (cc=147 and ll>=178 and ll<181) or (cc=148 and ll>=179 and ll<182) or (cc=149 and ll>=180 and ll<182) or (cc=150 and ll>=181 and ll<183) or (cc=151 and ll>=182 and ll<184) or (cc=152 and ll>=183 and ll<185) or (cc=153 and ll=185) or (cc=154 and ll>=185 and ll<187) or (cc=155 and ll>=186 and ll<188) or (cc=156 and ll=187) or (cc=157 and ll>=188 and ll<190) or (cc=158 and ll>=189 and ll<191) or (cc=159 and ll=190) or (cc=160 and ll=191) or (cc=161 and ll=192) or (cc=162 and ll=192)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0000")) then
	if ((cc=121 and ll>=158 and ll<161) or (cc=122 and ll>=153 and ll<162) or (cc=123 and ll>=154 and ll<163) or (cc=124 and ll>=155 and ll<165) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=157 and ll<165) or (cc=127 and ll>=158 and ll<166) or (cc=128 and ll>=160 and ll<167) or (cc=129 and ll>=161 and ll<168) or (cc=130 and ll>=162 and ll<169) or (cc=131 and ll>=163 and ll<171) or (cc=132 and ll>=164 and ll<172) or (cc=133 and ll>=167 and ll<173) or (cc=134 and ll>=168 and ll<174) or (cc=135 and ll>=169 and ll<175) or (cc=136 and ll>=170 and ll<176) or (cc=137 and ll>=171 and ll<177) or (cc=138 and ll>=172 and ll<179) or (cc=139 and ll>=173 and ll<180) or (cc=140 and ll>=175 and ll<181) or (cc=141 and ll>=176 and ll<182) or (cc=142 and ll>=178 and ll<183) or (cc=143 and ll>=179 and ll<184) or (cc=144 and ll>=181 and ll<186) or (cc=145 and ll>=182 and ll<186) or (cc=146 and ll>=183 and ll<185) or (cc=147 and ll>=184 and ll<186) or (cc=148 and ll>=185 and ll<188) or (cc=149 and ll>=186 and ll<189) or (cc=150 and ll>=187 and ll<190) or (cc=151 and ll>=189 and ll<191) or (cc=152 and ll=191) or (cc=153 and ll=192) or (cc=154 and ll>=193 and ll<195) or (cc=155 and ll>=194 and ll<196) or (cc=156 and ll>=195 and ll<197) or (cc=157 and ll>=196 and ll<198) or (cc=158 and ll>=197 and ll<199) or (cc=159 and ll=199) or (cc=160 and ll=200)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0001")) then
	if ((cc=121 and ll>=157 and ll<161) or (cc=122 and ll>=154 and ll<162) or (cc=123 and ll>=153 and ll<164) or (cc=124 and ll>=155 and ll<165) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=158 and ll<166) or (cc=127 and ll>=159 and ll<167) or (cc=128 and ll>=160 and ll<168) or (cc=129 and ll>=162 and ll<170) or (cc=130 and ll>=163 and ll<171) or (cc=131 and ll>=165 and ll<173) or (cc=132 and ll>=166 and ll<174) or (cc=133 and ll>=169 and ll<176) or (cc=134 and ll>=170 and ll<177) or (cc=135 and ll>=171 and ll<178) or (cc=136 and ll>=173 and ll<180) or (cc=137 and ll>=174 and ll<181) or (cc=138 and ll>=176 and ll<183) or (cc=139 and ll>=177 and ll<184) or (cc=140 and ll>=179 and ll<185) or (cc=141 and ll>=181 and ll<187) or (cc=142 and ll>=183 and ll<188) or (cc=143 and ll>=184 and ll<190) or (cc=144 and ll>=186 and ll<189) or (cc=145 and ll>=187 and ll<190) or (cc=146 and ll>=188 and ll<192) or (cc=147 and ll>=190 and ll<193) or (cc=148 and ll>=191 and ll<194) or (cc=149 and ll>=193 and ll<196) or (cc=150 and ll=196) or (cc=151 and ll>=197 and ll<199) or (cc=152 and ll=199) or (cc=153 and ll>=200 and ll<202) or (cc=154 and ll=202) or (cc=155 and ll>=203 and ll<205) or (cc=156 and ll=205) or (cc=157 and ll>=206 and ll<208)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0010")) then
	if ((cc=121 and ll>=156 and ll<160) or (cc=122 and ll>=154 and ll<161) or (cc=123 and ll>=152 and ll<163) or (cc=124 and ll>=154 and ll<165) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=157 and ll<166) or (cc=127 and ll>=159 and ll<168) or (cc=128 and ll>=161 and ll<170) or (cc=129 and ll>=162 and ll<171) or (cc=130 and ll>=164 and ll<173) or (cc=131 and ll>=166 and ll<175) or (cc=132 and ll>=169 and ll<176) or (cc=133 and ll>=171 and ll<178) or (cc=134 and ll>=173 and ll<181) or (cc=135 and ll>=175 and ll<182) or (cc=136 and ll>=177 and ll<184) or (cc=137 and ll>=179 and ll<186) or (cc=138 and ll>=180 and ll<188) or (cc=139 and ll>=182 and ll<189) or (cc=140 and ll>=185 and ll<191) or (cc=141 and ll>=187 and ll<193) or (cc=142 and ll>=189 and ll<194) or (cc=143 and ll>=191 and ll<194) or (cc=144 and ll>=192 and ll<196) or (cc=145 and ll>=194 and ll<198) or (cc=146 and ll>=196 and ll<199) or (cc=147 and ll>=197 and ll<201) or (cc=148 and ll>=201 and ll<203) or (cc=149 and ll=203) or (cc=150 and ll>=204 and ll<206) or (cc=151 and ll>=206 and ll<208) or (cc=152 and ll>=208 and ll<210) or (cc=153 and ll>=209 and ll<212) or (cc=154 and ll>=211 and ll<214) or (cc=155 and ll=213)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0011")) then
	if ((cc=121 and ll=157) or (cc=122 and ll>=154 and ll<161) or (cc=123 and ll>=152 and ll<163) or (cc=124 and ll>=153 and ll<165) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=157 and ll<167) or (cc=127 and ll>=159 and ll<169) or (cc=128 and ll>=162 and ll<171) or (cc=129 and ll>=164 and ll<173) or (cc=130 and ll>=166 and ll<176) or (cc=131 and ll>=168 and ll<178) or (cc=132 and ll>=172 and ll<180) or (cc=133 and ll>=174 and ll<182) or (cc=134 and ll>=176 and ll<185) or (cc=135 and ll>=179 and ll<187) or (cc=136 and ll>=181 and ll<189) or (cc=137 and ll>=183 and ll<191) or (cc=138 and ll>=185 and ll<193) or (cc=139 and ll>=189 and ll<196) or (cc=140 and ll>=191 and ll<197) or (cc=141 and ll>=193 and ll<197) or (cc=142 and ll>=196 and ll<200) or (cc=143 and ll>=198 and ll<202) or (cc=144 and ll>=200 and ll<204) or (cc=145 and ll>=202 and ll<206) or (cc=146 and ll>=206 and ll<208) or (cc=147 and ll>=208 and ll<211) or (cc=148 and ll>=210 and ll<213) or (cc=149 and ll>=213 and ll<215) or (cc=150 and ll>=215 and ll<217) or (cc=151 and ll>=216 and ll<219) or (cc=152 and ll=219)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0100")) then
	if ((cc=121 and ll>=156 and ll<158) or (cc=122 and ll>=155 and ll<160) or (cc=123 and ll>=152 and ll<163) or (cc=124 and ll>=152 and ll<166) or (cc=125 and ll>=154 and ll<165) or (cc=126 and ll>=157 and ll<168) or (cc=127 and ll>=159 and ll<171) or (cc=128 and ll>=162 and ll<173) or (cc=129 and ll>=165 and ll<176) or (cc=130 and ll>=168 and ll<179) or (cc=131 and ll>=172 and ll<182) or (cc=132 and ll>=175 and ll<185) or (cc=133 and ll>=177 and ll<187) or (cc=134 and ll>=181 and ll<190) or (cc=135 and ll>=183 and ll<193) or (cc=136 and ll>=185 and ll<195) or (cc=137 and ll>=190 and ll<199) or (cc=138 and ll>=193 and ll<200) or (cc=139 and ll>=196 and ll<201) or (cc=140 and ll>=198 and ll<203) or (cc=141 and ll>=201 and ll<205) or (cc=142 and ll>=204 and ll<209) or (cc=143 and ll>=206 and ll<211) or (cc=144 and ll>=211 and ll<214) or (cc=145 and ll>=214 and ll<217) or (cc=146 and ll>=217 and ll<219) or (cc=147 and ll>=219 and ll<222) or (cc=148 and ll>=222 and ll<225) or (cc=149 and ll=225)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0101")) then
	if ((cc=121 and ll=155) or (cc=122 and ll>=154 and ll<160) or (cc=123 and ll>=153 and ll<163) or (cc=124 and ll>=152 and ll<166) or (cc=125 and ll>=152 and ll<166) or (cc=126 and ll>=156 and ll<170) or (cc=127 and ll>=159 and ll<173) or (cc=128 and ll>=163 and ll<177) or (cc=129 and ll>=166 and ll<180) or (cc=130 and ll>=170 and ll<184) or (cc=131 and ll>=175 and ll<187) or (cc=132 and ll>=179 and ll<191) or (cc=133 and ll>=182 and ll<194) or (cc=134 and ll>=186 and ll<197) or (cc=135 and ll>=189 and ll<201) or (cc=136 and ll>=195 and ll<203) or (cc=137 and ll>=198 and ll<203) or (cc=138 and ll>=202 and ll<207) or (cc=139 and ll>=205 and ll<210) or (cc=140 and ll>=208 and ll<214) or (cc=141 and ll>=214 and ll<217) or (cc=142 and ll>=217 and ll<221) or (cc=143 and ll>=221 and ll<224) or (cc=144 and ll>=224 and ll<228) or (cc=145 and ll>=227 and ll<230)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0110")) then
	if ((cc=122 and ll>=154 and ll<159) or (cc=123 and ll>=153 and ll<164) or (cc=124 and ll>=152 and ll<165) or (cc=125 and ll>=151 and ll<167) or (cc=126 and ll>=155 and ll<172) or (cc=127 and ll>=160 and ll<176) or (cc=128 and ll>=164 and ll<181) or (cc=129 and ll>=169 and ll<186) or (cc=130 and ll>=176 and ll<190) or (cc=131 and ll>=180 and ll<195) or (cc=132 and ll>=185 and ll<199) or (cc=133 and ll>=189 and ll<203) or (cc=134 and ll>=196 and ll<205) or (cc=135 and ll>=201 and ll<208) or (cc=136 and ll>=205 and ll<212) or (cc=137 and ll>=209 and ll<217) or (cc=138 and ll>=217 and ll<220) or (cc=139 and ll>=220 and ll<225) or (cc=140 and ll>=225 and ll<229) or (cc=141 and ll>=229 and ll<234)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="0111")) then
	if ((cc=122 and ll>=154 and ll<158) or (cc=123 and ll>=153 and ll<164) or (cc=124 and ll>=152 and ll<165) or (cc=125 and ll>=151 and ll<170) or (cc=126 and ll>=154 and ll<176) or (cc=127 and ll>=160 and ll<183) or (cc=128 and ll>=166 and ll<188) or (cc=129 and ll>=172 and ll<194) or (cc=130 and ll>=181 and ll<201) or (cc=131 and ll>=188 and ll<206) or (cc=132 and ll>=194 and ll<207) or (cc=133 and ll>=203 and ll<212) or (cc=134 and ll>=209 and ll<218) or (cc=135 and ll>=215 and ll<225) or (cc=136 and ll>=225 and ll<230) or (cc=137 and ll>=230 and ll<237)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="1000")) then
	if ((cc=122 and ll>=153 and ll<156) or (cc=123 and ll>=153 and ll<165) or (cc=124 and ll>=152 and ll<165) or (cc=125 and ll>=152 and ll<175) or (cc=126 and ll>=152 and ll<184) or (cc=127 and ll>=160 and ll<193) or (cc=128 and ll>=169 and ll<202) or (cc=129 and ll>=183 and ll<207) or (cc=130 and ll>=193 and ll<212) or (cc=131 and ll>=207 and ll<221) or (cc=132 and ll>=216 and ll<230) or (cc=133 and ll>=230 and ll<239)) then grbp<="001";
	end if;

elsif ((PT2 ="0010" and PT3 ="1001")) then
	if ((cc=123 and ll>=152 and ll<164) or (cc=124 and ll>=152 and ll<170) or (cc=125 and ll>=152 and ll<188) or (cc=126 and ll>=152 and ll<207) or (cc=127 and ll>=161 and ll<208) or (cc=128 and ll>=188 and ll<226) or (cc=129 and ll>=216 and ll<241)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0000")) then
	if ((cc=123 and ll>=152 and ll<164) or (cc=124 and ll>=152 and ll<208) or (cc=125 and ll>=152 and ll<241) or (cc=126 and ll>=152 and ll<219) or (cc=127 and ll>=161 and ll<175)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0001")) then
	if ((cc=121 and ll>=230 and ll<241) or (cc=122 and ll>=190 and ll<230) or (cc=123 and ll>=152 and ll<219) or (cc=124 and ll>=152 and ll<200) or (cc=125 and ll>=152 and ll<190) or (cc=126 and ll>=152 and ll<175) or (cc=127 and ll>=152 and ll<160)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0010")) then
	if ((cc=117 and ll>=232 and ll<239) or (cc=118 and ll>=223 and ll<232) or (cc=119 and ll>=204 and ll<223) or (cc=120 and ll>=194 and ll<218) or (cc=121 and ll>=184 and ll<208) or (cc=122 and ll>=174 and ll<198) or (cc=123 and ll>=155 and ll<194) or (cc=124 and ll>=151 and ll<185) or (cc=125 and ll>=152 and ll<175) or (cc=126 and ll>=152 and ll<170) or (cc=127 and ll>=153 and ll<161)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0011")) then
	if ((cc=113 and ll>=232 and ll<237) or (cc=114 and ll>=226 and ll<232) or (cc=115 and ll>=220 and ll<226) or (cc=116 and ll>=213 and ll<220) or (cc=117 and ll>=200 and ll<217) or (cc=118 and ll>=195 and ll<211) or (cc=119 and ll>=188 and ll<204) or (cc=120 and ll>=182 and ll<198) or (cc=121 and ll>=176 and ll<195) or (cc=122 and ll>=170 and ll<189) or (cc=123 and ll>=157 and ll<183) or (cc=124 and ll>=151 and ll<177) or (cc=125 and ll>=152 and ll<173) or (cc=126 and ll>=152 and ll<168) or (cc=127 and ll>=153 and ll<161) or (cc=128 and ll=153)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0100")) then
	if ((cc=109 and ll>=230 and ll<234) or (cc=110 and ll>=226 and ll<231) or (cc=111 and ll>=221 and ll<226) or (cc=112 and ll>=217 and ll<221) or (cc=113 and ll>=212 and ll<217) or (cc=114 and ll>=208 and ll<214) or (cc=115 and ll>=199 and ll<211) or (cc=116 and ll>=194 and ll<206) or (cc=117 and ll>=189 and ll<202) or (cc=118 and ll>=185 and ll<197) or (cc=119 and ll>=180 and ll<195) or (cc=120 and ll>=176 and ll<190) or (cc=121 and ll>=171 and ll<186) or (cc=122 and ll>=167 and ll<181) or (cc=123 and ll>=157 and ll<176) or (cc=124 and ll>=153 and ll<175) or (cc=125 and ll>=151 and ll<170) or (cc=126 and ll>=152 and ll<166) or (cc=127 and ll>=153 and ll<161) or (cc=128 and ll>=153 and ll<157)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0101")) then
	if ((cc=105 and ll=229) or (cc=106 and ll>=225 and ll<229) or (cc=107 and ll>=222 and ll<225) or (cc=108 and ll>=218 and ll<222) or (cc=109 and ll>=215 and ll<218) or (cc=110 and ll>=211 and ll<215) or (cc=111 and ll>=208 and ll<212) or (cc=112 and ll>=200 and ll<210) or (cc=113 and ll>=196 and ll<207) or (cc=114 and ll>=193 and ll<203) or (cc=115 and ll>=189 and ll<199) or (cc=116 and ll>=186 and ll<195) or (cc=117 and ll>=182 and ll<193) or (cc=118 and ll>=179 and ll<191) or (cc=119 and ll>=175 and ll<187) or (cc=120 and ll>=172 and ll<184) or (cc=121 and ll>=169 and ll<180) or (cc=122 and ll>=165 and ll<177) or (cc=123 and ll>=158 and ll<175) or (cc=124 and ll>=155 and ll<172) or (cc=125 and ll>=151 and ll<169) or (cc=126 and ll>=152 and ll<165) or (cc=127 and ll>=153 and ll<162) or (cc=128 and ll>=154 and ll<158)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0110")) then
	if ((cc=102 and ll>=222 and ll<226) or (cc=103 and ll>=220 and ll<223) or (cc=104 and ll>=218 and ll<220) or (cc=105 and ll>=214 and ll<218) or (cc=106 and ll>=212 and ll<215) or (cc=107 and ll>=209 and ll<212) or (cc=108 and ll>=206 and ll<209) or (cc=109 and ll>=203 and ll<208) or (cc=110 and ll>=197 and ll<205) or (cc=111 and ll>=195 and ll<202) or (cc=112 and ll>=191 and ll<200) or (cc=113 and ll>=189 and ll<197) or (cc=114 and ll>=186 and ll<194) or (cc=115 and ll>=183 and ll<192) or (cc=116 and ll>=181 and ll<191) or (cc=117 and ll>=177 and ll<187) or (cc=118 and ll>=175 and ll<185) or (cc=119 and ll>=173 and ll<182) or (cc=120 and ll>=169 and ll<179) or (cc=121 and ll>=167 and ll<177) or (cc=122 and ll>=164 and ll<174) or (cc=123 and ll>=158 and ll<172) or (cc=124 and ll>=155 and ll<170) or (cc=125 and ll>=152 and ll<167) or (cc=126 and ll>=151 and ll<164) or (cc=127 and ll>=152 and ll<162) or (cc=128 and ll>=154 and ll<159) or (cc=129 and ll=155)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="0111")) then
	if ((cc=98 and ll=220) or (cc=99 and ll>=217 and ll<220) or (cc=100 and ll>=215 and ll<218) or (cc=101 and ll>=213 and ll<215) or (cc=102 and ll>=211 and ll<213) or (cc=103 and ll>=208 and ll<211) or (cc=104 and ll>=206 and ll<209) or (cc=105 and ll>=204 and ll<206) or (cc=106 and ll>=202 and ll<205) or (cc=107 and ll>=200 and ll<203) or (cc=108 and ll>=197 and ll<201) or (cc=109 and ll>=192 and ll<199) or (cc=110 and ll>=190 and ll<197) or (cc=111 and ll>=188 and ll<194) or (cc=112 and ll>=186 and ll<192) or (cc=113 and ll>=183 and ll<190) or (cc=114 and ll>=181 and ll<189) or (cc=115 and ll>=179 and ll<187) or (cc=116 and ll>=177 and ll<185) or (cc=117 and ll>=174 and ll<182) or (cc=118 and ll>=172 and ll<180) or (cc=119 and ll>=170 and ll<178) or (cc=120 and ll>=168 and ll<176) or (cc=121 and ll>=165 and ll<174) or (cc=122 and ll>=163 and ll<173) or (cc=123 and ll>=158 and ll<170) or (cc=124 and ll>=156 and ll<168) or (cc=125 and ll>=154 and ll<166) or (cc=126 and ll>=151 and ll<164) or (cc=127 and ll>=153 and ll<162) or (cc=128 and ll>=154 and ll<159) or (cc=129 and ll=156)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="1000")) then
	if ((cc=95 and ll=214) or (cc=96 and ll>=212 and ll<214) or (cc=97 and ll>=210 and ll<212) or (cc=98 and ll>=208 and ll<211) or (cc=99 and ll>=206 and ll<209) or (cc=100 and ll>=205 and ll<207) or (cc=101 and ll>=203 and ll<205) or (cc=102 and ll>=201 and ll<203) or (cc=103 and ll=200) or (cc=104 and ll>=198 and ll<201) or (cc=105 and ll>=196 and ll<199) or (cc=106 and ll>=194 and ll<197) or (cc=107 and ll>=189 and ll<195) or (cc=108 and ll>=187 and ll<194) or (cc=109 and ll>=186 and ll<192) or (cc=110 and ll>=184 and ll<190) or (cc=111 and ll>=182 and ll<189) or (cc=112 and ll>=180 and ll<187) or (cc=113 and ll>=179 and ll<186) or (cc=114 and ll>=177 and ll<184) or (cc=115 and ll>=175 and ll<183) or (cc=116 and ll>=173 and ll<181) or (cc=117 and ll>=171 and ll<179) or (cc=118 and ll>=169 and ll<177) or (cc=119 and ll>=168 and ll<175) or (cc=120 and ll>=166 and ll<173) or (cc=121 and ll>=164 and ll<173) or (cc=122 and ll>=162 and ll<171) or (cc=123 and ll>=158 and ll<169) or (cc=124 and ll>=156 and ll<167) or (cc=125 and ll>=154 and ll<166) or (cc=126 and ll>=152 and ll<164) or (cc=127 and ll>=152 and ll<162) or (cc=128 and ll>=155 and ll<160) or (cc=129 and ll>=156 and ll<159)) then grbp<="001";
	end if;

elsif ((PT2 ="0011" and PT3 ="1001")) then
	if ((cc=93 and ll=207) or (cc=94 and ll>=205 and ll<207) or (cc=95 and ll=204) or (cc=96 and ll>=202 and ll<204) or (cc=97 and ll=201) or (cc=98 and ll>=199 and ll<201) or (cc=99 and ll=198) or (cc=100 and ll>=196 and ll<198) or (cc=101 and ll=195) or (cc=102 and ll>=193 and ll<196) or (cc=103 and ll>=192 and ll<195) or (cc=104 and ll>=190 and ll<194) or (cc=105 and ll>=186 and ll<192) or (cc=106 and ll>=185 and ll<191) or (cc=107 and ll>=183 and ll<189) or (cc=108 and ll>=182 and ll<188) or (cc=109 and ll>=180 and ll<186) or (cc=110 and ll>=179 and ll<185) or (cc=111 and ll>=177 and ll<184) or (cc=112 and ll>=176 and ll<183) or (cc=113 and ll>=175 and ll<182) or (cc=114 and ll>=173 and ll<180) or (cc=115 and ll>=172 and ll<179) or (cc=116 and ll>=170 and ll<177) or (cc=117 and ll>=169 and ll<176) or (cc=118 and ll>=167 and ll<174) or (cc=119 and ll>=166 and ll<173) or (cc=120 and ll>=164 and ll<172) or (cc=121 and ll>=163 and ll<171) or (cc=122 and ll>=161 and ll<169) or (cc=123 and ll>=157 and ll<168) or (cc=124 and ll>=156 and ll<166) or (cc=125 and ll>=154 and ll<165) or (cc=126 and ll>=153 and ll<163) or (cc=127 and ll>=152 and ll<162) or (cc=128 and ll>=154 and ll<160) or (cc=129 and ll>=156 and ll<159)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0000")) then
	if ((cc=90 and ll=200) or (cc=91 and ll>=199 and ll<201) or (cc=92 and ll>=198 and ll<200) or (cc=93 and ll>=197 and ll<199) or (cc=94 and ll=196) or (cc=95 and ll=195) or (cc=96 and ll>=193 and ll<195) or (cc=97 and ll>=192 and ll<194) or (cc=98 and ll>=191 and ll<193) or (cc=99 and ll>=190 and ll<192) or (cc=100 and ll>=189 and ll<191) or (cc=101 and ll>=188 and ll<191) or (cc=102 and ll>=187 and ll<189) or (cc=103 and ll>=185 and ll<188) or (cc=104 and ll>=182 and ll<187) or (cc=105 and ll>=180 and ll<186) or (cc=106 and ll>=179 and ll<185) or (cc=107 and ll>=178 and ll<184) or (cc=108 and ll>=177 and ll<182) or (cc=109 and ll>=176 and ll<181) or (cc=110 and ll>=175 and ll<181) or (cc=111 and ll>=174 and ll<180) or (cc=112 and ll>=172 and ll<179) or (cc=113 and ll>=171 and ll<178) or (cc=114 and ll>=170 and ll<176) or (cc=115 and ll>=169 and ll<175) or (cc=116 and ll>=168 and ll<174) or (cc=117 and ll>=167 and ll<173) or (cc=118 and ll>=165 and ll<172) or (cc=119 and ll>=164 and ll<171) or (cc=120 and ll>=163 and ll<171) or (cc=121 and ll>=162 and ll<170) or (cc=122 and ll>=161 and ll<168) or (cc=123 and ll>=158 and ll<167) or (cc=124 and ll>=156 and ll<166) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=154 and ll<164) or (cc=127 and ll>=153 and ll<163) or (cc=128 and ll>=154 and ll<161) or (cc=129 and ll>=157 and ll<160)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0001")) then
	if ((cc=89 and ll>=192 and ll<194) or (cc=90 and ll>=191 and ll<193) or (cc=91 and ll>=190 and ll<192) or (cc=92 and ll=190) or (cc=93 and ll=189) or (cc=94 and ll>=187 and ll<189) or (cc=95 and ll=187) or (cc=96 and ll=186) or (cc=97 and ll=185) or (cc=98 and ll>=184 and ll<186) or (cc=99 and ll>=183 and ll<186) or (cc=100 and ll>=182 and ll<185) or (cc=101 and ll>=181 and ll<184) or (cc=102 and ll>=181 and ll<183) or (cc=103 and ll>=177 and ll<182) or (cc=104 and ll>=177 and ll<181) or (cc=105 and ll>=175 and ll<180) or (cc=106 and ll>=175 and ll<180) or (cc=107 and ll>=174 and ll<179) or (cc=108 and ll>=173 and ll<177) or (cc=109 and ll>=172 and ll<178) or (cc=110 and ll>=171 and ll<177) or (cc=111 and ll>=170 and ll<176) or (cc=112 and ll>=169 and ll<175) or (cc=113 and ll>=168 and ll<174) or (cc=114 and ll>=168 and ll<173) or (cc=115 and ll>=166 and ll<172) or (cc=116 and ll>=166 and ll<171) or (cc=117 and ll>=165 and ll<171) or (cc=118 and ll>=164 and ll<170) or (cc=119 and ll>=163 and ll<169) or (cc=120 and ll>=162 and ll<169) or (cc=121 and ll>=161 and ll<168) or (cc=122 and ll>=160 and ll<167) or (cc=123 and ll>=157 and ll<166) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=156 and ll<165) or (cc=126 and ll>=154 and ll<164) or (cc=127 and ll>=153 and ll<163) or (cc=128 and ll>=153 and ll<162) or (cc=129 and ll>=157 and ll<161)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0010")) then
	if ((cc=87 and ll=185) or (cc=88 and ll=184) or (cc=89 and ll>=183 and ll<185) or (cc=90 and ll=183) or (cc=91 and ll>=182 and ll<184) or (cc=92 and ll=182) or (cc=93 and ll=181) or (cc=94 and ll>=180 and ll<182) or (cc=95 and ll=180) or (cc=96 and ll=179) or (cc=97 and ll>=178 and ll<180) or (cc=98 and ll>=178 and ll<180) or (cc=99 and ll>=177 and ll<179) or (cc=100 and ll>=176 and ll<179) or (cc=101 and ll>=176 and ll<178) or (cc=102 and ll>=173 and ll<177) or (cc=103 and ll>=172 and ll<177) or (cc=104 and ll>=172 and ll<176) or (cc=105 and ll>=171 and ll<175) or (cc=106 and ll>=170 and ll<175) or (cc=107 and ll>=170 and ll<174) or (cc=108 and ll>=169 and ll<174) or (cc=109 and ll>=168 and ll<174) or (cc=110 and ll>=167 and ll<173) or (cc=111 and ll>=167 and ll<173) or (cc=112 and ll>=166 and ll<172) or (cc=113 and ll>=166 and ll<171) or (cc=114 and ll>=165 and ll<170) or (cc=115 and ll>=164 and ll<170) or (cc=116 and ll>=164 and ll<169) or (cc=117 and ll>=163 and ll<169) or (cc=118 and ll>=162 and ll<168) or (cc=119 and ll>=162 and ll<168) or (cc=120 and ll>=161 and ll<168) or (cc=121 and ll>=160 and ll<167) or (cc=122 and ll>=160 and ll<166) or (cc=123 and ll>=157 and ll<166) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=155 and ll<164) or (cc=127 and ll>=154 and ll<163) or (cc=128 and ll>=154 and ll<162) or (cc=129 and ll>=157 and ll<162)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0011")) then
	if ((cc=86 and ll=177) or (cc=87 and ll>=176 and ll<178) or (cc=88 and ll=176) or (cc=89 and ll>=175 and ll<177) or (cc=90 and ll=175) or (cc=91 and ll=175) or (cc=92 and ll=174) or (cc=93 and ll=174) or (cc=94 and ll>=173 and ll<175) or (cc=95 and ll=173) or (cc=96 and ll>=172 and ll<174) or (cc=97 and ll>=172 and ll<174) or (cc=98 and ll>=172 and ll<174) or (cc=99 and ll>=171 and ll<173) or (cc=100 and ll>=171 and ll<173) or (cc=101 and ll>=170 and ll<173) or (cc=102 and ll>=168 and ll<172) or (cc=103 and ll>=167 and ll<172) or (cc=104 and ll>=167 and ll<171) or (cc=105 and ll>=167 and ll<171) or (cc=106 and ll>=166 and ll<170) or (cc=107 and ll>=166 and ll<170) or (cc=108 and ll>=165 and ll<171) or (cc=109 and ll>=165 and ll<170) or (cc=110 and ll>=164 and ll<170) or (cc=111 and ll>=164 and ll<169) or (cc=112 and ll>=164 and ll<169) or (cc=113 and ll>=163 and ll<168) or (cc=114 and ll>=163 and ll<168) or (cc=115 and ll>=162 and ll<167) or (cc=116 and ll>=162 and ll<167) or (cc=117 and ll>=161 and ll<167) or (cc=118 and ll>=161 and ll<167) or (cc=119 and ll>=160 and ll<167) or (cc=120 and ll>=160 and ll<166) or (cc=121 and ll>=160 and ll<166) or (cc=122 and ll>=159 and ll<165) or (cc=123 and ll>=157 and ll<165) or (cc=124 and ll>=156 and ll<165) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=155 and ll<164) or (cc=127 and ll>=155 and ll<163) or (cc=128 and ll>=154 and ll<163) or (cc=129 and ll>=156 and ll<162)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0100")) then
	if ((cc=85 and ll=169) or (cc=86 and ll>=168 and ll<170) or (cc=87 and ll=168) or (cc=88 and ll=168) or (cc=89 and ll=168) or (cc=90 and ll=168) or (cc=91 and ll=167) or (cc=92 and ll=167) or (cc=93 and ll=167) or (cc=94 and ll=167) or (cc=95 and ll=167) or (cc=96 and ll>=166 and ll<168) or (cc=97 and ll>=166 and ll<168) or (cc=98 and ll>=166 and ll<168) or (cc=99 and ll>=166 and ll<168) or (cc=100 and ll>=165 and ll<168) or (cc=101 and ll>=165 and ll<167) or (cc=102 and ll>=163 and ll<167) or (cc=103 and ll>=163 and ll<167) or (cc=104 and ll>=163 and ll<167) or (cc=105 and ll>=162 and ll<166) or (cc=106 and ll>=162 and ll<166) or (cc=107 and ll>=162 and ll<167) or (cc=108 and ll>=162 and ll<167) or (cc=109 and ll>=161 and ll<167) or (cc=110 and ll>=161 and ll<166) or (cc=111 and ll>=161 and ll<166) or (cc=112 and ll>=161 and ll<166) or (cc=113 and ll>=161 and ll<166) or (cc=114 and ll>=160 and ll<165) or (cc=115 and ll>=160 and ll<165) or (cc=116 and ll>=160 and ll<165) or (cc=117 and ll>=160 and ll<165) or (cc=118 and ll>=159 and ll<166) or (cc=119 and ll>=159 and ll<165) or (cc=120 and ll>=159 and ll<165) or (cc=121 and ll>=159 and ll<165) or (cc=122 and ll>=159 and ll<165) or (cc=123 and ll>=156 and ll<165) or (cc=124 and ll>=156 and ll<164) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=156 and ll<164) or (cc=127 and ll>=155 and ll<164) or (cc=128 and ll>=155 and ll<163) or (cc=129 and ll>=155 and ll<163)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0101")) then
	if ((cc=85 and ll=160) or (cc=86 and ll=160) or (cc=87 and ll=160) or (cc=88 and ll=160) or (cc=89 and ll=160) or (cc=90 and ll=160) or (cc=91 and ll=160) or (cc=92 and ll=160) or (cc=93 and ll=160) or (cc=94 and ll=160) or (cc=95 and ll=160) or (cc=96 and ll>=160 and ll<162) or (cc=97 and ll>=160 and ll<162) or (cc=98 and ll>=160 and ll<162) or (cc=99 and ll>=160 and ll<162) or (cc=100 and ll>=160 and ll<162) or (cc=101 and ll>=158 and ll<162) or (cc=102 and ll>=158 and ll<162) or (cc=103 and ll>=158 and ll<162) or (cc=104 and ll>=158 and ll<162) or (cc=105 and ll>=158 and ll<162) or (cc=106 and ll>=158 and ll<162) or (cc=107 and ll>=158 and ll<163) or (cc=108 and ll>=158 and ll<163) or (cc=109 and ll>=158 and ll<163) or (cc=110 and ll>=158 and ll<163) or (cc=111 and ll>=158 and ll<163) or (cc=112 and ll>=158 and ll<163) or (cc=113 and ll>=158 and ll<163) or (cc=114 and ll>=158 and ll<163) or (cc=115 and ll>=158 and ll<163) or (cc=116 and ll>=158 and ll<163) or (cc=117 and ll>=158 and ll<163) or (cc=118 and ll>=158 and ll<164) or (cc=119 and ll>=158 and ll<164) or (cc=120 and ll>=158 and ll<164) or (cc=121 and ll>=158 and ll<164) or (cc=122 and ll>=158 and ll<164) or (cc=123 and ll>=156 and ll<164) or (cc=124 and ll>=156 and ll<164) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=156 and ll<164) or (cc=127 and ll>=156 and ll<164) or (cc=128 and ll>=156 and ll<164) or (cc=129 and ll>=156 and ll<164)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0110")) then
	if ((cc=85 and ll=152) or (cc=86 and ll=152) or (cc=87 and ll=152) or (cc=88 and ll>=152 and ll<154) or (cc=89 and ll=153) or (cc=90 and ll=153) or (cc=91 and ll=153) or (cc=92 and ll=153) or (cc=93 and ll>=153 and ll<155) or (cc=94 and ll=154) or (cc=95 and ll=154) or (cc=96 and ll>=154 and ll<156) or (cc=97 and ll>=154 and ll<156) or (cc=98 and ll>=154 and ll<157) or (cc=99 and ll>=155 and ll<157) or (cc=100 and ll>=155 and ll<157) or (cc=101 and ll>=155 and ll<157) or (cc=102 and ll>=153 and ll<157) or (cc=103 and ll>=153 and ll<158) or (cc=104 and ll>=154 and ll<158) or (cc=105 and ll>=154 and ll<158) or (cc=106 and ll>=154 and ll<158) or (cc=107 and ll>=154 and ll<159) or (cc=108 and ll>=154 and ll<160) or (cc=109 and ll>=155 and ll<160) or (cc=110 and ll>=155 and ll<160) or (cc=111 and ll>=155 and ll<160) or (cc=112 and ll>=155 and ll<160) or (cc=113 and ll>=155 and ll<161) or (cc=114 and ll>=156 and ll<161) or (cc=115 and ll>=156 and ll<161) or (cc=116 and ll>=156 and ll<161) or (cc=117 and ll>=156 and ll<161) or (cc=118 and ll>=157 and ll<163) or (cc=119 and ll>=157 and ll<163) or (cc=120 and ll>=157 and ll<163) or (cc=121 and ll>=157 and ll<163) or (cc=122 and ll>=157 and ll<163) or (cc=123 and ll>=158 and ll<164) or (cc=124 and ll>=156 and ll<164) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=156 and ll<164) or (cc=127 and ll>=156 and ll<164) or (cc=128 and ll>=157 and ll<165) or (cc=129 and ll>=157 and ll<165)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="0111")) then
	if ((cc=86 and ll=144) or (cc=87 and ll=144) or (cc=88 and ll=145) or (cc=89 and ll=145) or (cc=90 and ll>=145 and ll<147) or (cc=91 and ll=146) or (cc=92 and ll=146) or (cc=93 and ll=147) or (cc=94 and ll=147) or (cc=95 and ll>=147 and ll<149) or (cc=96 and ll=148) or (cc=97 and ll>=148 and ll<151) or (cc=98 and ll>=149 and ll<151) or (cc=99 and ll>=149 and ll<151) or (cc=100 and ll>=149 and ll<152) or (cc=101 and ll>=150 and ll<152) or (cc=102 and ll>=148 and ll<153) or (cc=103 and ll>=149 and ll<153) or (cc=104 and ll>=149 and ll<153) or (cc=105 and ll>=149 and ll<154) or (cc=106 and ll>=150 and ll<154) or (cc=107 and ll>=150 and ll<156) or (cc=108 and ll>=151 and ll<156) or (cc=109 and ll>=151 and ll<156) or (cc=110 and ll>=152 and ll<157) or (cc=111 and ll>=152 and ll<157) or (cc=112 and ll>=153 and ll<158) or (cc=113 and ll>=153 and ll<158) or (cc=114 and ll>=153 and ll<158) or (cc=115 and ll>=154 and ll<159) or (cc=116 and ll>=154 and ll<159) or (cc=117 and ll>=155 and ll<160) or (cc=118 and ll>=155 and ll<161) or (cc=119 and ll>=155 and ll<162) or (cc=120 and ll>=156 and ll<162) or (cc=121 and ll>=156 and ll<163) or (cc=122 and ll>=157 and ll<163) or (cc=123 and ll>=157 and ll<163) or (cc=124 and ll>=155 and ll<164) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=157 and ll<165) or (cc=128 and ll>=157 and ll<165) or (cc=129 and ll>=158 and ll<166)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="1000")) then
	if ((cc=87 and ll=136) or (cc=88 and ll>=136 and ll<138) or (cc=89 and ll=137) or (cc=90 and ll>=137 and ll<139) or (cc=91 and ll=138) or (cc=92 and ll=139) or (cc=93 and ll>=139 and ll<141) or (cc=94 and ll=140) or (cc=95 and ll>=140 and ll<142) or (cc=96 and ll>=141 and ll<143) or (cc=97 and ll>=142 and ll<144) or (cc=98 and ll>=143 and ll<145) or (cc=99 and ll>=143 and ll<145) or (cc=100 and ll>=144 and ll<146) or (cc=101 and ll>=144 and ll<147) or (cc=102 and ll>=145 and ll<148) or (cc=103 and ll>=144 and ll<148) or (cc=104 and ll>=144 and ll<149) or (cc=105 and ll>=145 and ll<149) or (cc=106 and ll>=146 and ll<150) or (cc=107 and ll>=146 and ll<151) or (cc=108 and ll>=147 and ll<152) or (cc=109 and ll>=147 and ll<153) or (cc=110 and ll>=148 and ll<154) or (cc=111 and ll>=149 and ll<154) or (cc=112 and ll>=150 and ll<155) or (cc=113 and ll>=150 and ll<156) or (cc=114 and ll>=151 and ll<156) or (cc=115 and ll>=151 and ll<157) or (cc=116 and ll>=152 and ll<157) or (cc=117 and ll>=153 and ll<158) or (cc=118 and ll>=153 and ll<160) or (cc=119 and ll>=154 and ll<161) or (cc=120 and ll>=154 and ll<161) or (cc=121 and ll>=155 and ll<162) or (cc=122 and ll>=156 and ll<162) or (cc=123 and ll>=157 and ll<163) or (cc=124 and ll>=155 and ll<164) or (cc=125 and ll>=156 and ll<164) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=157 and ll<166) or (cc=128 and ll>=157 and ll<166) or (cc=129 and ll>=158 and ll<165)) then grbp<="001";
	end if;

elsif ((PT2 ="0100" and PT3 ="1001")) then
	if ((cc=88 and ll=128) or (cc=89 and ll>=128 and ll<130) or (cc=90 and ll=129) or (cc=91 and ll=130) or (cc=92 and ll=131) or (cc=93 and ll>=131 and ll<133) or (cc=94 and ll=133) or (cc=95 and ll>=133 and ll<135) or (cc=96 and ll>=134 and ll<136) or (cc=97 and ll=135) or (cc=98 and ll>=136 and ll<139) or (cc=99 and ll>=137 and ll<139) or (cc=100 and ll>=138 and ll<140) or (cc=101 and ll>=139 and ll<141) or (cc=102 and ll>=139 and ll<142) or (cc=103 and ll>=140 and ll<143) or (cc=104 and ll>=139 and ll<144) or (cc=105 and ll>=140 and ll<145) or (cc=106 and ll>=141 and ll<146) or (cc=107 and ll>=142 and ll<147) or (cc=108 and ll>=142 and ll<148) or (cc=109 and ll>=144 and ll<150) or (cc=110 and ll>=144 and ll<150) or (cc=111 and ll>=145 and ll<151) or (cc=112 and ll>=146 and ll<152) or (cc=113 and ll>=147 and ll<153) or (cc=114 and ll>=148 and ll<154) or (cc=115 and ll>=149 and ll<155) or (cc=116 and ll>=150 and ll<156) or (cc=117 and ll>=151 and ll<156) or (cc=118 and ll>=151 and ll<159) or (cc=119 and ll>=152 and ll<159) or (cc=120 and ll>=153 and ll<160) or (cc=121 and ll>=154 and ll<161) or (cc=122 and ll>=155 and ll<162) or (cc=123 and ll>=156 and ll<163) or (cc=124 and ll>=155 and ll<164) or (cc=125 and ll>=156 and ll<165) or (cc=126 and ll>=156 and ll<165) or (cc=127 and ll>=157 and ll<166) or (cc=128 and ll>=158 and ll<167) or (cc=129 and ll>=159 and ll<164)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0000")) then
	if ((cc=90 and ll=120) or (cc=91 and ll=121) or (cc=92 and ll>=122 and ll<124) or (cc=93 and ll>=123 and ll<125) or (cc=94 and ll>=124 and ll<126) or (cc=95 and ll>=125 and ll<127) or (cc=96 and ll=127) or (cc=97 and ll=128) or (cc=98 and ll=129) or (cc=99 and ll>=130 and ll<132) or (cc=100 and ll>=131 and ll<134) or (cc=101 and ll>=132 and ll<135) or (cc=102 and ll>=133 and ll<136) or (cc=103 and ll>=135 and ll<138) or (cc=104 and ll>=136 and ll<139) or (cc=105 and ll>=135 and ll<140) or (cc=106 and ll>=135 and ll<141) or (cc=107 and ll>=137 and ll<142) or (cc=108 and ll>=138 and ll<143) or (cc=109 and ll>=139 and ll<145) or (cc=110 and ll>=140 and ll<146) or (cc=111 and ll>=141 and ll<148) or (cc=112 and ll>=142 and ll<149) or (cc=113 and ll>=144 and ll<150) or (cc=114 and ll>=145 and ll<151) or (cc=115 and ll>=146 and ll<152) or (cc=116 and ll>=147 and ll<153) or (cc=117 and ll>=148 and ll<154) or (cc=118 and ll>=149 and ll<157) or (cc=119 and ll>=150 and ll<158) or (cc=120 and ll>=152 and ll<159) or (cc=121 and ll>=153 and ll<160) or (cc=122 and ll>=154 and ll<161) or (cc=123 and ll>=155 and ll<163) or (cc=124 and ll>=156 and ll<164) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=156 and ll<166) or (cc=127 and ll>=158 and ll<167) or (cc=128 and ll>=159 and ll<168) or (cc=129 and ll>=160 and ll<163)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0001")) then
	if ((cc=93 and ll>=113 and ll<115) or (cc=94 and ll>=115 and ll<117) or (cc=95 and ll>=116 and ll<118) or (cc=96 and ll>=118 and ll<120) or (cc=97 and ll>=119 and ll<121) or (cc=98 and ll=121) or (cc=99 and ll>=122 and ll<124) or (cc=100 and ll=124) or (cc=101 and ll>=125 and ll<128) or (cc=102 and ll>=127 and ll<130) or (cc=103 and ll>=128 and ll<131) or (cc=104 and ll>=130 and ll<133) or (cc=105 and ll>=131 and ll<134) or (cc=106 and ll>=132 and ll<136) or (cc=107 and ll>=131 and ll<137) or (cc=108 and ll>=133 and ll<138) or (cc=109 and ll>=134 and ll<140) or (cc=110 and ll>=136 and ll<142) or (cc=111 and ll>=137 and ll<144) or (cc=112 and ll>=139 and ll<145) or (cc=113 and ll>=140 and ll<147) or (cc=114 and ll>=141 and ll<148) or (cc=115 and ll>=143 and ll<150) or (cc=116 and ll>=144 and ll<151) or (cc=117 and ll>=146 and ll<152) or (cc=118 and ll>=147 and ll<155) or (cc=119 and ll>=148 and ll<156) or (cc=120 and ll>=150 and ll<158) or (cc=121 and ll>=151 and ll<159) or (cc=122 and ll>=153 and ll<161) or (cc=123 and ll>=154 and ll<162) or (cc=124 and ll>=155 and ll<163) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=156 and ll<166) or (cc=127 and ll>=157 and ll<168) or (cc=128 and ll>=159 and ll<167) or (cc=129 and ll>=160 and ll<164)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0010")) then
	if ((cc=95 and ll=107) or (cc=96 and ll>=107 and ll<110) or (cc=97 and ll>=109 and ll<112) or (cc=98 and ll>=111 and ll<113) or (cc=99 and ll>=113 and ll<115) or (cc=100 and ll>=115 and ll<117) or (cc=101 and ll>=117 and ll<119) or (cc=102 and ll=119) or (cc=103 and ll>=120 and ll<124) or (cc=104 and ll>=122 and ll<125) or (cc=105 and ll>=124 and ll<127) or (cc=106 and ll>=125 and ll<129) or (cc=107 and ll>=127 and ll<130) or (cc=108 and ll>=127 and ll<132) or (cc=109 and ll>=128 and ll<134) or (cc=110 and ll>=130 and ll<136) or (cc=111 and ll>=132 and ll<139) or (cc=112 and ll>=134 and ll<141) or (cc=113 and ll>=135 and ll<143) or (cc=114 and ll>=137 and ll<145) or (cc=115 and ll>=139 and ll<147) or (cc=116 and ll>=141 and ll<148) or (cc=117 and ll>=143 and ll<150) or (cc=118 and ll>=145 and ll<152) or (cc=119 and ll>=146 and ll<155) or (cc=120 and ll>=148 and ll<157) or (cc=121 and ll>=150 and ll<159) or (cc=122 and ll>=151 and ll<160) or (cc=123 and ll>=153 and ll<162) or (cc=124 and ll>=155 and ll<164) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=156 and ll<167) or (cc=127 and ll>=158 and ll<169) or (cc=128 and ll>=160 and ll<167) or (cc=129 and ll>=161 and ll<165)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0011")) then
	if ((cc=98 and ll>=101 and ll<103) or (cc=99 and ll>=102 and ll<105) or (cc=100 and ll>=104 and ll<107) or (cc=101 and ll>=107 and ll<109) or (cc=102 and ll>=109 and ll<111) or (cc=103 and ll>=111 and ll<114) or (cc=104 and ll>=113 and ll<116) or (cc=105 and ll>=116 and ll<119) or (cc=106 and ll>=117 and ll<122) or (cc=107 and ll>=119 and ll<124) or (cc=108 and ll>=122 and ll<126) or (cc=109 and ll>=124 and ll<128) or (cc=110 and ll>=124 and ll<130) or (cc=111 and ll>=125 and ll<132) or (cc=112 and ll>=128 and ll<136) or (cc=113 and ll>=130 and ll<138) or (cc=114 and ll>=132 and ll<140) or (cc=115 and ll>=134 and ll<142) or (cc=116 and ll>=136 and ll<145) or (cc=117 and ll>=139 and ll<147) or (cc=118 and ll>=141 and ll<149) or (cc=119 and ll>=143 and ll<153) or (cc=120 and ll>=145 and ll<155) or (cc=121 and ll>=148 and ll<157) or (cc=122 and ll>=150 and ll<159) or (cc=123 and ll>=152 and ll<162) or (cc=124 and ll>=154 and ll<164) or (cc=125 and ll>=155 and ll<166) or (cc=126 and ll>=156 and ll<168) or (cc=127 and ll>=158 and ll<169) or (cc=128 and ll>=160 and ll<167) or (cc=129 and ll>=162 and ll<164)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0100")) then
	if ((cc=101 and ll=95) or (cc=102 and ll>=96 and ll<99) or (cc=103 and ll>=99 and ll<102) or (cc=104 and ll>=102 and ll<105) or (cc=105 and ll>=104 and ll<108) or (cc=106 and ll>=108 and ll<110) or (cc=107 and ll>=110 and ll<115) or (cc=108 and ll>=112 and ll<117) or (cc=109 and ll>=116 and ll<120) or (cc=110 and ll>=118 and ll<123) or (cc=111 and ll>=120 and ll<125) or (cc=112 and ll>=121 and ll<129) or (cc=113 and ll>=123 and ll<131) or (cc=114 and ll>=126 and ll<136) or (cc=115 and ll>=128 and ll<138) or (cc=116 and ll>=131 and ll<140) or (cc=117 and ll>=134 and ll<144) or (cc=118 and ll>=136 and ll<146) or (cc=119 and ll>=139 and ll<149) or (cc=120 and ll>=142 and ll<153) or (cc=121 and ll>=145 and ll<156) or (cc=122 and ll>=148 and ll<159) or (cc=123 and ll>=150 and ll<162) or (cc=124 and ll>=153 and ll<164) or (cc=125 and ll>=156 and ll<167) or (cc=126 and ll>=155 and ll<169) or (cc=127 and ll>=158 and ll<169) or (cc=128 and ll>=161 and ll<166) or (cc=129 and ll>=163 and ll<165)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0101")) then
	if ((cc=105 and ll>=91 and ll<94) or (cc=106 and ll>=93 and ll<97) or (cc=107 and ll>=97 and ll<101) or (cc=108 and ll>=100 and ll<104) or (cc=109 and ll>=104 and ll<107) or (cc=110 and ll>=107 and ll<113) or (cc=111 and ll>=111 and ll<117) or (cc=112 and ll>=114 and ll<120) or (cc=113 and ll>=118 and ll<123) or (cc=114 and ll>=118 and ll<127) or (cc=115 and ll>=120 and ll<132) or (cc=116 and ll>=124 and ll<135) or (cc=117 and ll>=127 and ll<139) or (cc=118 and ll>=130 and ll<142) or (cc=119 and ll>=134 and ll<146) or (cc=120 and ll>=137 and ll<151) or (cc=121 and ll>=141 and ll<155) or (cc=122 and ll>=144 and ll<158) or (cc=123 and ll>=148 and ll<162) or (cc=124 and ll>=151 and ll<165) or (cc=125 and ll>=155 and ll<169) or (cc=126 and ll>=155 and ll<169) or (cc=127 and ll>=158 and ll<168) or (cc=128 and ll>=161 and ll<167) or (cc=129 and ll=165)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0110")) then
	if ((cc=109 and ll>=87 and ll<92) or (cc=110 and ll>=92 and ll<96) or (cc=111 and ll>=96 and ll<101) or (cc=112 and ll>=101 and ll<105) or (cc=113 and ll>=105 and ll<112) or (cc=114 and ll>=110 and ll<117) or (cc=115 and ll>=114 and ll<120) or (cc=116 and ll>=116 and ll<125) or (cc=117 and ll>=118 and ll<132) or (cc=118 and ll>=123 and ll<136) or (cc=119 and ll>=126 and ll<141) or (cc=120 and ll>=131 and ll<145) or (cc=121 and ll>=135 and ll<152) or (cc=122 and ll>=140 and ll<157) or (cc=123 and ll>=145 and ll<161) or (cc=124 and ll>=149 and ll<166) or (cc=125 and ll>=154 and ll<170) or (cc=126 and ll>=156 and ll<169) or (cc=127 and ll>=157 and ll<168) or (cc=128 and ll>=162 and ll<167)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="0111")) then
	if ((cc=112 and ll=84) or (cc=113 and ll>=85 and ll<91) or (cc=114 and ll>=91 and ll<96) or (cc=115 and ll>=96 and ll<106) or (cc=116 and ll>=103 and ll<112) or (cc=117 and ll>=109 and ll<119) or (cc=118 and ll>=115 and ll<127) or (cc=119 and ll>=115 and ll<133) or (cc=120 and ll>=120 and ll<140) or (cc=121 and ll>=127 and ll<149) or (cc=122 and ll>=133 and ll<155) or (cc=123 and ll>=138 and ll<161) or (cc=124 and ll>=145 and ll<167) or (cc=125 and ll>=151 and ll<170) or (cc=126 and ll>=156 and ll<169) or (cc=127 and ll>=157 and ll<168) or (cc=128 and ll>=163 and ll<167)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="1000")) then
	if ((cc=117 and ll>=82 and ll<92) or (cc=118 and ll>=92 and ll<106) or (cc=119 and ll>=100 and ll<114) or (cc=120 and ll>=110 and ll<128) or (cc=121 and ll>=114 and ll<138) or (cc=122 and ll>=119 and ll<152) or (cc=123 and ll>=128 and ll<161) or (cc=124 and ll>=137 and ll<169) or (cc=125 and ll>=147 and ll<169) or (cc=126 and ll>=156 and ll<169) or (cc=127 and ll>=156 and ll<168) or (cc=128 and ll>=165 and ll<168)) then grbp<="001";
	end if;

elsif ((PT2 ="0101" and PT3 ="1001")) then
	if ((cc=121 and ll>=80 and ll<106) or (cc=122 and ll>=96 and ll<133) or (cc=123 and ll>=113 and ll<160) or (cc=124 and ll>=115 and ll<169) or (cc=125 and ll>=133 and ll<169) or (cc=126 and ll>=151 and ll<169) or (cc=127 and ll>=157 and ll<169)) then grbp<="001";
	end if;


end if;
if ((PT4 ="0000" and PT5 ="0000")) then
	if ((cc=122 and ll>=156 and ll<160) or (cc=123 and ll>=112 and ll<173) or (cc=124 and ll>=68 and ll<173) or (cc=125 and ll>=46 and ll<173) or (cc=126 and ll>=79 and ll<173) or (cc=127 and ll>=123 and ll<173) or (cc=128 and ll>=167 and ll<173)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0001")) then
	if ((cc=122 and ll>=160 and ll<173) or (cc=123 and ll>=151 and ll<173) or (cc=124 and ll>=134 and ll<173) or (cc=125 and ll>=122 and ll<173) or (cc=126 and ll>=112 and ll<173) or (cc=127 and ll>=93 and ll<174) or (cc=128 and ll>=83 and ll<171) or (cc=129 and ll>=68 and ll<132) or (cc=130 and ll>=55 and ll<93) or (cc=131 and ll>=47 and ll<55)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0010")) then
	if ((cc=121 and ll>=170 and ll<172) or (cc=122 and ll>=160 and ll<172) or (cc=123 and ll>=155 and ll<173) or (cc=124 and ll>=145 and ll<173) or (cc=125 and ll>=137 and ll<173) or (cc=126 and ll>=132 and ll<174) or (cc=127 and ll>=122 and ll<174) or (cc=128 and ll>=112 and ll<156) or (cc=129 and ll>=108 and ll<147) or (cc=130 and ll>=99 and ll<137) or (cc=131 and ll>=91 and ll<128) or (cc=132 and ll>=84 and ll<109) or (cc=133 and ll>=75 and ll<99) or (cc=134 and ll>=70 and ll<90) or (cc=135 and ll>=61 and ll<70) or (cc=136 and ll>=51 and ll<61) or (cc=137 and ll>=48 and ll<51)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0011")) then
	if ((cc=121 and ll>=166 and ll<171) or (cc=122 and ll>=159 and ll<172) or (cc=123 and ll>=155 and ll<172) or (cc=124 and ll>=150 and ll<173) or (cc=125 and ll>=144 and ll<174) or (cc=126 and ll>=138 and ll<174) or (cc=127 and ll>=134 and ll<170) or (cc=128 and ll>=129 and ll<158) or (cc=129 and ll>=123 and ll<152) or (cc=130 and ll>=116 and ll<146) or (cc=131 and ll>=113 and ll<139) or (cc=132 and ll>=108 and ll<134) or (cc=133 and ll>=101 and ll<127) or (cc=134 and ll>=95 and ll<114) or (cc=135 and ll>=92 and ll<108) or (cc=136 and ll>=86 and ll<102) or (cc=137 and ll>=80 and ll<96) or (cc=138 and ll>=74 and ll<89) or (cc=139 and ll>=71 and ll<77) or (cc=140 and ll>=65 and ll<71) or (cc=141 and ll>=58 and ll<65) or (cc=142 and ll>=52 and ll<58) or (cc=143 and ll=52)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0100")) then
	if ((cc=120 and ll>=168 and ll<170) or (cc=121 and ll>=163 and ll<171) or (cc=122 and ll>=160 and ll<172) or (cc=123 and ll>=155 and ll<173) or (cc=124 and ll>=153 and ll<174) or (cc=125 and ll>=148 and ll<174) or (cc=126 and ll>=144 and ll<173) or (cc=127 and ll>=139 and ll<164) or (cc=128 and ll>=135 and ll<159) or (cc=129 and ll>=133 and ll<154) or (cc=130 and ll>=129 and ll<150) or (cc=131 and ll>=124 and ll<145) or (cc=132 and ll>=119 and ll<141) or (cc=133 and ll>=115 and ll<136) or (cc=134 and ll>=113 and ll<132) or (cc=135 and ll>=108 and ll<122) or (cc=136 and ll>=103 and ll<118) or (cc=137 and ll>=99 and ll<113) or (cc=138 and ll>=95 and ll<109) or (cc=139 and ll>=93 and ll<104) or (cc=140 and ll>=88 and ll<100) or (cc=141 and ll>=84 and ll<95) or (cc=142 and ll>=79 and ll<91) or (cc=143 and ll>=75 and ll<81) or (cc=144 and ll>=72 and ll<77) or (cc=145 and ll>=68 and ll<72) or (cc=146 and ll>=63 and ll<68) or (cc=147 and ll>=59 and ll<63) or (cc=148 and ll>=56 and ll<59)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0101")) then
	if ((cc=120 and ll>=166 and ll<169) or (cc=121 and ll>=163 and ll<170) or (cc=122 and ll>=159 and ll<171) or (cc=123 and ll>=156 and ll<172) or (cc=124 and ll>=154 and ll<173) or (cc=125 and ll>=151 and ll<174) or (cc=126 and ll>=148 and ll<171) or (cc=127 and ll>=144 and ll<163) or (cc=128 and ll>=140 and ll<160) or (cc=129 and ll>=136 and ll<156) or (cc=130 and ll>=135 and ll<153) or (cc=131 and ll>=132 and ll<149) or (cc=132 and ll>=128 and ll<146) or (cc=133 and ll>=125 and ll<142) or (cc=134 and ll>=121 and ll<139) or (cc=135 and ll>=118 and ll<135) or (cc=136 and ll>=117 and ll<132) or (cc=137 and ll>=113 and ll<125) or (cc=138 and ll>=110 and ll<121) or (cc=139 and ll>=106 and ll<118) or (cc=140 and ll>=103 and ll<114) or (cc=141 and ll>=99 and ll<111) or (cc=142 and ll>=98 and ll<107) or (cc=143 and ll>=94 and ll<104) or (cc=144 and ll>=91 and ll<100) or (cc=145 and ll>=87 and ll<97) or (cc=146 and ll>=83 and ll<94) or (cc=147 and ll>=80 and ll<86) or (cc=148 and ll>=79 and ll<82) or (cc=149 and ll>=75 and ll<79) or (cc=150 and ll>=72 and ll<75) or (cc=151 and ll>=68 and ll<72) or (cc=152 and ll>=65 and ll<68) or (cc=153 and ll>=61 and ll<65)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0110")) then
	if ((cc=119 and ll=167) or (cc=120 and ll>=164 and ll<169) or (cc=121 and ll>=162 and ll<171) or (cc=122 and ll>=159 and ll<172) or (cc=123 and ll>=156 and ll<173) or (cc=124 and ll>=154 and ll<174) or (cc=125 and ll>=152 and ll<172) or (cc=126 and ll>=150 and ll<166) or (cc=127 and ll>=146 and ll<163) or (cc=128 and ll>=144 and ll<160) or (cc=129 and ll>=141 and ll<158) or (cc=130 and ll>=138 and ll<155) or (cc=131 and ll>=137 and ll<152) or (cc=132 and ll>=135 and ll<150) or (cc=133 and ll>=132 and ll<146) or (cc=134 and ll>=129 and ll<144) or (cc=135 and ll>=127 and ll<141) or (cc=136 and ll>=123 and ll<138) or (cc=137 and ll>=121 and ll<136) or (cc=138 and ll>=119 and ll<130) or (cc=139 and ll>=117 and ll<127) or (cc=140 and ll>=114 and ll<124) or (cc=141 and ll>=111 and ll<121) or (cc=142 and ll>=109 and ll<118) or (cc=143 and ll>=106 and ll<116) or (cc=144 and ll>=103 and ll<113) or (cc=145 and ll>=102 and ll<110) or (cc=146 and ll>=99 and ll<107) or (cc=147 and ll>=96 and ll<105) or (cc=148 and ll>=94 and ll<102) or (cc=149 and ll>=91 and ll<99) or (cc=150 and ll>=88 and ll<97) or (cc=151 and ll>=86 and ll<91) or (cc=152 and ll>=85 and ll<87) or (cc=153 and ll>=81 and ll<85) or (cc=154 and ll>=79 and ll<82) or (cc=155 and ll>=76 and ll<79) or (cc=156 and ll>=73 and ll<76) or (cc=157 and ll>=71 and ll<74) or (cc=158 and ll>=68 and ll<71)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="0111")) then
	if ((cc=119 and ll>=165 and ll<167) or (cc=120 and ll>=163 and ll<169) or (cc=121 and ll>=160 and ll<170) or (cc=122 and ll>=158 and ll<173) or (cc=123 and ll>=156 and ll<174) or (cc=124 and ll>=154 and ll<173) or (cc=125 and ll>=154 and ll<171) or (cc=126 and ll>=151 and ll<165) or (cc=127 and ll>=149 and ll<163) or (cc=128 and ll>=147 and ll<161) or (cc=129 and ll>=145 and ll<158) or (cc=130 and ll>=142 and ll<156) or (cc=131 and ll>=140 and ll<154) or (cc=132 and ll>=138 and ll<152) or (cc=133 and ll>=137 and ll<150) or (cc=134 and ll>=135 and ll<147) or (cc=135 and ll>=133 and ll<146) or (cc=136 and ll>=130 and ll<144) or (cc=137 and ll>=128 and ll<141) or (cc=138 and ll>=126 and ll<139) or (cc=139 and ll>=124 and ll<137) or (cc=140 and ll>=122 and ll<131) or (cc=141 and ll>=121 and ll<129) or (cc=142 and ll>=118 and ll<127) or (cc=143 and ll>=116 and ll<124) or (cc=144 and ll>=114 and ll<122) or (cc=145 and ll>=112 and ll<120) or (cc=146 and ll>=110 and ll<118) or (cc=147 and ll>=107 and ll<115) or (cc=148 and ll>=106 and ll<113) or (cc=149 and ll>=104 and ll<111) or (cc=150 and ll>=102 and ll<109) or (cc=151 and ll>=100 and ll<107) or (cc=152 and ll>=98 and ll<104) or (cc=153 and ll>=95 and ll<102) or (cc=154 and ll>=93 and ll<97) or (cc=155 and ll>=91 and ll<95) or (cc=156 and ll>=90 and ll<93) or (cc=157 and ll>=88 and ll<90) or (cc=158 and ll>=86 and ll<88) or (cc=159 and ll>=83 and ll<86) or (cc=160 and ll>=81 and ll<84) or (cc=161 and ll>=79 and ll<81) or (cc=162 and ll>=77 and ll<79) or (cc=163 and ll>=75 and ll<77)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="1000")) then
	if ((cc=119 and ll>=164 and ll<166) or (cc=120 and ll>=162 and ll<168) or (cc=121 and ll>=160 and ll<171) or (cc=122 and ll>=158 and ll<172) or (cc=123 and ll>=156 and ll<173) or (cc=124 and ll>=154 and ll<171) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=152 and ll<165) or (cc=127 and ll>=150 and ll<163) or (cc=128 and ll>=148 and ll<161) or (cc=129 and ll>=147 and ll<160) or (cc=130 and ll>=145 and ll<158) or (cc=131 and ll>=143 and ll<156) or (cc=132 and ll>=142 and ll<155) or (cc=133 and ll>=140 and ll<153) or (cc=134 and ll>=139 and ll<151) or (cc=135 and ll>=137 and ll<149) or (cc=136 and ll>=136 and ll<147) or (cc=137 and ll>=134 and ll<145) or (cc=138 and ll>=132 and ll<143) or (cc=139 and ll>=130 and ll<142) or (cc=140 and ll>=128 and ll<140) or (cc=141 and ll>=126 and ll<136) or (cc=142 and ll>=126 and ll<134) or (cc=143 and ll>=124 and ll<132) or (cc=144 and ll>=122 and ll<130) or (cc=145 and ll>=120 and ll<128) or (cc=146 and ll>=119 and ll<126) or (cc=147 and ll>=117 and ll<124) or (cc=148 and ll>=115 and ll<123) or (cc=149 and ll>=114 and ll<121) or (cc=150 and ll>=112 and ll<119) or (cc=151 and ll>=111 and ll<118) or (cc=152 and ll>=109 and ll<116) or (cc=153 and ll>=108 and ll<114) or (cc=154 and ll>=106 and ll<112) or (cc=155 and ll>=104 and ll<110) or (cc=156 and ll>=102 and ll<108) or (cc=157 and ll>=100 and ll<104) or (cc=158 and ll>=98 and ll<102) or (cc=159 and ll>=98 and ll<100) or (cc=160 and ll>=96 and ll<98) or (cc=161 and ll>=94 and ll<97) or (cc=162 and ll>=92 and ll<95) or (cc=163 and ll>=91 and ll<93) or (cc=164 and ll>=89 and ll<91) or (cc=165 and ll>=87 and ll<89) or (cc=166 and ll=86) or (cc=167 and ll>=84 and ll<86)) then grbp<="101";
	end if;

elsif ((PT4 ="0000" and PT5 ="1001")) then
	if ((cc=119 and ll>=162 and ll<166) or (cc=120 and ll>=161 and ll<168) or (cc=121 and ll>=159 and ll<171) or (cc=122 and ll>=158 and ll<173) or (cc=123 and ll>=157 and ll<172) or (cc=124 and ll>=155 and ll<171) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=153 and ll<165) or (cc=127 and ll>=151 and ll<164) or (cc=128 and ll>=150 and ll<162) or (cc=129 and ll>=149 and ll<161) or (cc=130 and ll>=147 and ll<159) or (cc=131 and ll>=146 and ll<158) or (cc=132 and ll>=144 and ll<156) or (cc=133 and ll>=143 and ll<155) or (cc=134 and ll>=141 and ll<153) or (cc=135 and ll>=141 and ll<152) or (cc=136 and ll>=140 and ll<150) or (cc=137 and ll>=138 and ll<149) or (cc=138 and ll>=137 and ll<147) or (cc=139 and ll>=135 and ll<146) or (cc=140 and ll>=134 and ll<145) or (cc=141 and ll>=132 and ll<143) or (cc=142 and ll>=131 and ll<139) or (cc=143 and ll>=130 and ll<138) or (cc=144 and ll>=129 and ll<136) or (cc=145 and ll>=128 and ll<135) or (cc=146 and ll>=127 and ll<133) or (cc=147 and ll>=125 and ll<132) or (cc=148 and ll>=124 and ll<130) or (cc=149 and ll>=122 and ll<129) or (cc=150 and ll>=121 and ll<127) or (cc=151 and ll>=119 and ll<126) or (cc=152 and ll>=118 and ll<124) or (cc=153 and ll>=117 and ll<123) or (cc=154 and ll>=116 and ll<121) or (cc=155 and ll>=114 and ll<120) or (cc=156 and ll>=113 and ll<118) or (cc=157 and ll>=111 and ll<117) or (cc=158 and ll>=110 and ll<115) or (cc=159 and ll>=108 and ll<112) or (cc=160 and ll>=107 and ll<110) or (cc=161 and ll>=106 and ll<109) or (cc=162 and ll>=105 and ll<107) or (cc=163 and ll>=104 and ll<106) or (cc=164 and ll=103) or (cc=165 and ll>=101 and ll<103) or (cc=166 and ll=100) or (cc=167 and ll>=98 and ll<100) or (cc=168 and ll>=97 and ll<99) or (cc=169 and ll>=95 and ll<97) or (cc=170 and ll>=94 and ll<96) or (cc=171 and ll=93)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0000")) then
	if ((cc=119 and ll>=161 and ll<165) or (cc=120 and ll>=160 and ll<169) or (cc=121 and ll>=159 and ll<172) or (cc=122 and ll>=157 and ll<172) or (cc=123 and ll>=156 and ll<171) or (cc=124 and ll>=155 and ll<167) or (cc=125 and ll>=154 and ll<166) or (cc=126 and ll>=154 and ll<165) or (cc=127 and ll>=153 and ll<163) or (cc=128 and ll>=152 and ll<162) or (cc=129 and ll>=151 and ll<161) or (cc=130 and ll>=149 and ll<160) or (cc=131 and ll>=148 and ll<159) or (cc=132 and ll>=147 and ll<158) or (cc=133 and ll>=146 and ll<156) or (cc=134 and ll>=144 and ll<155) or (cc=135 and ll>=143 and ll<154) or (cc=136 and ll>=143 and ll<153) or (cc=137 and ll>=142 and ll<152) or (cc=138 and ll>=141 and ll<151) or (cc=139 and ll>=140 and ll<150) or (cc=140 and ll>=139 and ll<148) or (cc=141 and ll>=138 and ll<147) or (cc=142 and ll>=136 and ll<146) or (cc=143 and ll>=135 and ll<143) or (cc=144 and ll>=134 and ll<142) or (cc=145 and ll>=133 and ll<141) or (cc=146 and ll>=133 and ll<139) or (cc=147 and ll>=132 and ll<138) or (cc=148 and ll>=131 and ll<137) or (cc=149 and ll>=130 and ll<136) or (cc=150 and ll>=128 and ll<135) or (cc=151 and ll>=127 and ll<134) or (cc=152 and ll>=126 and ll<132) or (cc=153 and ll>=125 and ll<131) or (cc=154 and ll>=124 and ll<130) or (cc=155 and ll>=123 and ll<129) or (cc=156 and ll>=123 and ll<128) or (cc=157 and ll>=121 and ll<127) or (cc=158 and ll>=120 and ll<126) or (cc=159 and ll>=119 and ll<124) or (cc=160 and ll>=118 and ll<123) or (cc=161 and ll>=117 and ll<122) or (cc=162 and ll>=115 and ll<118) or (cc=163 and ll>=114 and ll<117) or (cc=164 and ll>=113 and ll<116) or (cc=165 and ll>=113 and ll<115) or (cc=166 and ll>=112 and ll<114) or (cc=167 and ll>=111 and ll<113) or (cc=168 and ll=110) or (cc=169 and ll=109) or (cc=170 and ll>=107 and ll<109) or (cc=171 and ll>=106 and ll<108) or (cc=172 and ll>=105 and ll<107) or (cc=173 and ll>=104 and ll<106) or (cc=174 and ll=103)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0001")) then
	if ((cc=119 and ll>=160 and ll<165) or (cc=120 and ll>=159 and ll<170) or (cc=121 and ll>=158 and ll<171) or (cc=122 and ll>=157 and ll<171) or (cc=123 and ll>=156 and ll<170) or (cc=124 and ll>=155 and ll<167) or (cc=125 and ll>=154 and ll<165) or (cc=126 and ll>=154 and ll<165) or (cc=127 and ll>=153 and ll<164) or (cc=128 and ll>=153 and ll<163) or (cc=129 and ll>=152 and ll<162) or (cc=130 and ll>=151 and ll<161) or (cc=131 and ll>=150 and ll<160) or (cc=132 and ll>=149 and ll<159) or (cc=133 and ll>=148 and ll<159) or (cc=134 and ll>=147 and ll<158) or (cc=135 and ll>=147 and ll<156) or (cc=136 and ll>=146 and ll<156) or (cc=137 and ll>=146 and ll<155) or (cc=138 and ll>=145 and ll<154) or (cc=139 and ll>=144 and ll<153) or (cc=140 and ll>=143 and ll<152) or (cc=141 and ll>=142 and ll<151) or (cc=142 and ll>=141 and ll<150) or (cc=143 and ll>=141 and ll<150) or (cc=144 and ll>=139 and ll<146) or (cc=145 and ll>=138 and ll<146) or (cc=146 and ll>=138 and ll<144) or (cc=147 and ll>=138 and ll<144) or (cc=148 and ll>=137 and ll<143) or (cc=149 and ll>=136 and ll<142) or (cc=150 and ll>=135 and ll<141) or (cc=151 and ll>=134 and ll<140) or (cc=152 and ll>=133 and ll<139) or (cc=153 and ll>=132 and ll<138) or (cc=154 and ll>=132 and ll<137) or (cc=155 and ll>=131 and ll<137) or (cc=156 and ll>=130 and ll<136) or (cc=157 and ll>=130 and ll<135) or (cc=158 and ll>=129 and ll<134) or (cc=159 and ll>=128 and ll<133) or (cc=160 and ll>=127 and ll<132) or (cc=161 and ll>=126 and ll<131) or (cc=162 and ll>=126 and ll<130) or (cc=163 and ll>=125 and ll<127) or (cc=164 and ll>=124 and ll<126) or (cc=165 and ll>=123 and ll<125) or (cc=166 and ll>=122 and ll<125) or (cc=167 and ll>=121 and ll<124) or (cc=168 and ll>=121 and ll<123) or (cc=169 and ll>=120 and ll<122) or (cc=170 and ll=120) or (cc=171 and ll=119) or (cc=172 and ll>=117 and ll<119) or (cc=173 and ll=117) or (cc=174 and ll=116) or (cc=175 and ll=115) or (cc=176 and ll>=114 and ll<116) or (cc=177 and ll>=113 and ll<115)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0010")) then
	if ((cc=119 and ll>=158 and ll<165) or (cc=120 and ll>=158 and ll<170) or (cc=121 and ll>=157 and ll<170) or (cc=122 and ll>=156 and ll<170) or (cc=123 and ll>=156 and ll<169) or (cc=124 and ll>=155 and ll<166) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=154 and ll<165) or (cc=127 and ll>=154 and ll<164) or (cc=128 and ll>=154 and ll<164) or (cc=129 and ll>=153 and ll<163) or (cc=130 and ll>=152 and ll<162) or (cc=131 and ll>=152 and ll<161) or (cc=132 and ll>=151 and ll<161) or (cc=133 and ll>=150 and ll<160) or (cc=134 and ll>=150 and ll<160) or (cc=135 and ll>=149 and ll<159) or (cc=136 and ll>=148 and ll<158) or (cc=137 and ll>=148 and ll<158) or (cc=138 and ll>=148 and ll<157) or (cc=139 and ll>=148 and ll<156) or (cc=140 and ll>=147 and ll<155) or (cc=141 and ll>=146 and ll<155) or (cc=142 and ll>=146 and ll<154) or (cc=143 and ll>=145 and ll<154) or (cc=144 and ll>=144 and ll<151) or (cc=145 and ll>=143 and ll<150) or (cc=146 and ll>=143 and ll<150) or (cc=147 and ll>=142 and ll<149) or (cc=148 and ll>=143 and ll<148) or (cc=149 and ll>=142 and ll<148) or (cc=150 and ll>=141 and ll<147) or (cc=151 and ll>=141 and ll<146) or (cc=152 and ll>=140 and ll<145) or (cc=153 and ll>=139 and ll<145) or (cc=154 and ll>=139 and ll<144) or (cc=155 and ll>=138 and ll<144) or (cc=156 and ll>=138 and ll<143) or (cc=157 and ll>=137 and ll<142) or (cc=158 and ll>=136 and ll<142) or (cc=159 and ll>=137 and ll<141) or (cc=160 and ll>=136 and ll<140) or (cc=161 and ll>=135 and ll<140) or (cc=162 and ll>=134 and ll<139) or (cc=163 and ll>=134 and ll<138) or (cc=164 and ll>=133 and ll<138) or (cc=165 and ll>=133 and ll<135) or (cc=166 and ll>=132 and ll<134) or (cc=167 and ll>=131 and ll<134) or (cc=168 and ll>=131 and ll<133) or (cc=169 and ll>=130 and ll<132) or (cc=170 and ll>=130 and ll<132) or (cc=171 and ll=130) or (cc=172 and ll>=129 and ll<131) or (cc=173 and ll>=128 and ll<130) or (cc=174 and ll=128) or (cc=175 and ll=127) or (cc=176 and ll>=126 and ll<128) or (cc=177 and ll=126) or (cc=178 and ll=125) or (cc=179 and ll=125)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0011")) then
	if ((cc=119 and ll>=157 and ll<165) or (cc=120 and ll>=157 and ll<169) or (cc=121 and ll>=157 and ll<169) or (cc=122 and ll>=156 and ll<169) or (cc=123 and ll>=156 and ll<166) or (cc=124 and ll>=155 and ll<166) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=154 and ll<165) or (cc=127 and ll>=155 and ll<164) or (cc=128 and ll>=154 and ll<164) or (cc=129 and ll>=154 and ll<163) or (cc=130 and ll>=154 and ll<163) or (cc=131 and ll>=153 and ll<163) or (cc=132 and ll>=153 and ll<162) or (cc=133 and ll>=152 and ll<162) or (cc=134 and ll>=152 and ll<161) or (cc=135 and ll>=151 and ll<161) or (cc=136 and ll>=151 and ll<160) or (cc=137 and ll>=151 and ll<160) or (cc=138 and ll>=151 and ll<160) or (cc=139 and ll>=151 and ll<159) or (cc=140 and ll>=150 and ll<159) or (cc=141 and ll>=150 and ll<158) or (cc=142 and ll>=150 and ll<158) or (cc=143 and ll>=149 and ll<158) or (cc=144 and ll>=149 and ll<157) or (cc=145 and ll>=148 and ll<155) or (cc=146 and ll>=148 and ll<154) or (cc=147 and ll>=147 and ll<154) or (cc=148 and ll>=147 and ll<153) or (cc=149 and ll>=148 and ll<153) or (cc=150 and ll>=147 and ll<152) or (cc=151 and ll>=147 and ll<152) or (cc=152 and ll>=146 and ll<152) or (cc=153 and ll>=146 and ll<151) or (cc=154 and ll>=145 and ll<151) or (cc=155 and ll>=145 and ll<150) or (cc=156 and ll>=145 and ll<150) or (cc=157 and ll>=144 and ll<149) or (cc=158 and ll>=144 and ll<149) or (cc=159 and ll>=143 and ll<148) or (cc=160 and ll>=144 and ll<148) or (cc=161 and ll>=143 and ll<148) or (cc=162 and ll>=143 and ll<147) or (cc=163 and ll>=143 and ll<147) or (cc=164 and ll>=142 and ll<146) or (cc=165 and ll>=142 and ll<146) or (cc=166 and ll>=141 and ll<144) or (cc=167 and ll>=141 and ll<143) or (cc=168 and ll>=140 and ll<143) or (cc=169 and ll>=140 and ll<142) or (cc=170 and ll>=140 and ll<142) or (cc=171 and ll=140) or (cc=172 and ll=140) or (cc=173 and ll=139) or (cc=174 and ll=139) or (cc=175 and ll>=138 and ll<140) or (cc=176 and ll=138) or (cc=177 and ll=138) or (cc=178 and ll=137) or (cc=179 and ll=137) or (cc=180 and ll=136) or (cc=181 and ll=136)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0100")) then
	if ((cc=119 and ll>=156 and ll<168) or (cc=120 and ll>=156 and ll<168) or (cc=121 and ll>=156 and ll<168) or (cc=122 and ll>=156 and ll<168) or (cc=123 and ll>=155 and ll<166) or (cc=124 and ll>=155 and ll<165) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=155 and ll<165) or (cc=127 and ll>=155 and ll<165) or (cc=128 and ll>=155 and ll<164) or (cc=129 and ll>=155 and ll<164) or (cc=130 and ll>=155 and ll<164) or (cc=131 and ll>=155 and ll<164) or (cc=132 and ll>=154 and ll<164) or (cc=133 and ll>=154 and ll<163) or (cc=134 and ll>=154 and ll<163) or (cc=135 and ll>=154 and ll<163) or (cc=136 and ll>=154 and ll<163) or (cc=137 and ll>=153 and ll<163) or (cc=138 and ll>=153 and ll<162) or (cc=139 and ll>=154 and ll<162) or (cc=140 and ll>=154 and ll<162) or (cc=141 and ll>=153 and ll<162) or (cc=142 and ll>=153 and ll<161) or (cc=143 and ll>=153 and ll<161) or (cc=144 and ll>=153 and ll<161) or (cc=145 and ll>=153 and ll<159) or (cc=146 and ll>=152 and ll<159) or (cc=147 and ll>=152 and ll<158) or (cc=148 and ll>=152 and ll<158) or (cc=149 and ll>=152 and ll<158) or (cc=150 and ll>=153 and ll<158) or (cc=151 and ll>=152 and ll<157) or (cc=152 and ll>=152 and ll<157) or (cc=153 and ll>=152 and ll<157) or (cc=154 and ll>=152 and ll<157) or (cc=155 and ll>=151 and ll<157) or (cc=156 and ll>=151 and ll<156) or (cc=157 and ll>=151 and ll<156) or (cc=158 and ll>=151 and ll<156) or (cc=159 and ll>=151 and ll<156) or (cc=160 and ll>=151 and ll<156) or (cc=161 and ll>=151 and ll<155) or (cc=162 and ll>=151 and ll<155) or (cc=163 and ll>=151 and ll<155) or (cc=164 and ll>=151 and ll<155) or (cc=165 and ll>=150 and ll<154) or (cc=166 and ll>=150 and ll<152) or (cc=167 and ll>=150 and ll<152) or (cc=168 and ll>=150 and ll<152) or (cc=169 and ll>=149 and ll<152) or (cc=170 and ll>=149 and ll<151) or (cc=171 and ll>=149 and ll<151) or (cc=172 and ll=150) or (cc=173 and ll=150) or (cc=174 and ll>=149 and ll<151) or (cc=175 and ll=149) or (cc=176 and ll=149) or (cc=177 and ll=149) or (cc=178 and ll=149) or (cc=179 and ll=148) or (cc=180 and ll=148) or (cc=181 and ll=148) or (cc=182 and ll=148)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0101")) then
	if ((cc=119 and ll>=155 and ll<167) or (cc=120 and ll>=155 and ll<167) or (cc=121 and ll>=155 and ll<167) or (cc=122 and ll>=155 and ll<167) or (cc=123 and ll>=155 and ll<165) or (cc=124 and ll>=155 and ll<165) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=155 and ll<165) or (cc=127 and ll>=155 and ll<165) or (cc=128 and ll>=156 and ll<165) or (cc=129 and ll>=156 and ll<165) or (cc=130 and ll>=156 and ll<165) or (cc=131 and ll>=156 and ll<165) or (cc=132 and ll>=156 and ll<165) or (cc=133 and ll>=156 and ll<165) or (cc=134 and ll>=156 and ll<165) or (cc=135 and ll>=156 and ll<165) or (cc=136 and ll>=156 and ll<165) or (cc=137 and ll>=156 and ll<165) or (cc=138 and ll>=156 and ll<165) or (cc=139 and ll>=157 and ll<165) or (cc=140 and ll>=157 and ll<165) or (cc=141 and ll>=157 and ll<165) or (cc=142 and ll>=157 and ll<165) or (cc=143 and ll>=157 and ll<165) or (cc=144 and ll>=157 and ll<165) or (cc=145 and ll>=157 and ll<163) or (cc=146 and ll>=157 and ll<163) or (cc=147 and ll>=157 and ll<163) or (cc=148 and ll>=157 and ll<163) or (cc=149 and ll>=157 and ll<163) or (cc=150 and ll>=158 and ll<163) or (cc=151 and ll>=158 and ll<163) or (cc=152 and ll>=158 and ll<163) or (cc=153 and ll>=158 and ll<163) or (cc=154 and ll>=158 and ll<163) or (cc=155 and ll>=158 and ll<163) or (cc=156 and ll>=158 and ll<163) or (cc=157 and ll>=158 and ll<163) or (cc=158 and ll>=158 and ll<163) or (cc=159 and ll>=158 and ll<163) or (cc=160 and ll>=158 and ll<163) or (cc=161 and ll>=159 and ll<163) or (cc=162 and ll>=159 and ll<163) or (cc=163 and ll>=159 and ll<163) or (cc=164 and ll>=159 and ll<163) or (cc=165 and ll>=159 and ll<163) or (cc=166 and ll>=159 and ll<163) or (cc=167 and ll>=159 and ll<161) or (cc=168 and ll>=159 and ll<161) or (cc=169 and ll>=159 and ll<161) or (cc=170 and ll>=159 and ll<161) or (cc=171 and ll>=159 and ll<161) or (cc=172 and ll=160) or (cc=173 and ll=160) or (cc=174 and ll=160) or (cc=175 and ll=160) or (cc=176 and ll=160) or (cc=177 and ll=160) or (cc=178 and ll=160) or (cc=179 and ll=160) or (cc=180 and ll=160) or (cc=181 and ll=160) or (cc=182 and ll=160)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0110")) then
	if ((cc=119 and ll>=154 and ll<166) or (cc=120 and ll>=154 and ll<166) or (cc=121 and ll>=154 and ll<166) or (cc=122 and ll>=154 and ll<164) or (cc=123 and ll>=155 and ll<165) or (cc=124 and ll>=155 and ll<165) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=155 and ll<165) or (cc=127 and ll>=155 and ll<165) or (cc=128 and ll>=157 and ll<166) or (cc=129 and ll>=157 and ll<166) or (cc=130 and ll>=157 and ll<166) or (cc=131 and ll>=157 and ll<166) or (cc=132 and ll>=157 and ll<167) or (cc=133 and ll>=158 and ll<167) or (cc=134 and ll>=158 and ll<167) or (cc=135 and ll>=158 and ll<167) or (cc=136 and ll>=158 and ll<167) or (cc=137 and ll>=158 and ll<168) or (cc=138 and ll>=159 and ll<168) or (cc=139 and ll>=160 and ll<168) or (cc=140 and ll>=160 and ll<168) or (cc=141 and ll>=160 and ll<168) or (cc=142 and ll>=160 and ll<169) or (cc=143 and ll>=161 and ll<169) or (cc=144 and ll>=161 and ll<167) or (cc=145 and ll>=161 and ll<167) or (cc=146 and ll>=161 and ll<167) or (cc=147 and ll>=161 and ll<168) or (cc=148 and ll>=162 and ll<168) or (cc=149 and ll>=162 and ll<168) or (cc=150 and ll>=163 and ll<168) or (cc=151 and ll>=163 and ll<168) or (cc=152 and ll>=164 and ll<169) or (cc=153 and ll>=164 and ll<169) or (cc=154 and ll>=164 and ll<169) or (cc=155 and ll>=164 and ll<169) or (cc=156 and ll>=164 and ll<169) or (cc=157 and ll>=165 and ll<170) or (cc=158 and ll>=165 and ll<170) or (cc=159 and ll>=165 and ll<170) or (cc=160 and ll>=165 and ll<170) or (cc=161 and ll>=166 and ll<170) or (cc=162 and ll>=167 and ll<171) or (cc=163 and ll>=167 and ll<171) or (cc=164 and ll>=167 and ll<171) or (cc=165 and ll>=167 and ll<171) or (cc=166 and ll>=167 and ll<169) or (cc=167 and ll>=168 and ll<170) or (cc=168 and ll>=168 and ll<170) or (cc=169 and ll>=168 and ll<170) or (cc=170 and ll>=168 and ll<170) or (cc=171 and ll>=168 and ll<170) or (cc=172 and ll=170) or (cc=173 and ll=170) or (cc=174 and ll=170) or (cc=175 and ll=170) or (cc=176 and ll>=170 and ll<172) or (cc=177 and ll=171) or (cc=178 and ll=171) or (cc=179 and ll=171) or (cc=180 and ll=171) or (cc=181 and ll>=171 and ll<173) or (cc=182 and ll=172)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="0111")) then
	if ((cc=119 and ll>=155 and ll<165) or (cc=120 and ll>=153 and ll<165) or (cc=121 and ll>=153 and ll<165) or (cc=122 and ll>=153 and ll<164) or (cc=123 and ll>=154 and ll<164) or (cc=124 and ll>=154 and ll<165) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=155 and ll<166) or (cc=127 and ll>=156 and ll<166) or (cc=128 and ll>=157 and ll<166) or (cc=129 and ll>=158 and ll<167) or (cc=130 and ll>=158 and ll<167) or (cc=131 and ll>=158 and ll<168) or (cc=132 and ll>=159 and ll<168) or (cc=133 and ll>=159 and ll<169) or (cc=134 and ll>=160 and ll<169) or (cc=135 and ll>=160 and ll<169) or (cc=136 and ll>=160 and ll<170) or (cc=137 and ll>=161 and ll<170) or (cc=138 and ll>=161 and ll<171) or (cc=139 and ll>=163 and ll<171) or (cc=140 and ll>=163 and ll<171) or (cc=141 and ll>=164 and ll<172) or (cc=142 and ll>=164 and ll<172) or (cc=143 and ll>=164 and ll<173) or (cc=144 and ll>=165 and ll<171) or (cc=145 and ll>=165 and ll<172) or (cc=146 and ll>=166 and ll<172) or (cc=147 and ll>=166 and ll<172) or (cc=148 and ll>=167 and ll<173) or (cc=149 and ll>=167 and ll<173) or (cc=150 and ll>=168 and ll<174) or (cc=151 and ll>=169 and ll<174) or (cc=152 and ll>=169 and ll<174) or (cc=153 and ll>=170 and ll<175) or (cc=154 and ll>=170 and ll<175) or (cc=155 and ll>=170 and ll<176) or (cc=156 and ll>=171 and ll<176) or (cc=157 and ll>=171 and ll<177) or (cc=158 and ll>=172 and ll<177) or (cc=159 and ll>=172 and ll<177) or (cc=160 and ll>=174 and ll<178) or (cc=161 and ll>=174 and ll<178) or (cc=162 and ll>=174 and ll<179) or (cc=163 and ll>=175 and ll<179) or (cc=164 and ll>=175 and ll<180) or (cc=165 and ll>=176 and ll<178) or (cc=166 and ll>=176 and ll<178) or (cc=167 and ll>=176 and ll<179) or (cc=168 and ll>=177 and ll<179) or (cc=169 and ll>=177 and ll<179) or (cc=170 and ll>=178 and ll<180) or (cc=171 and ll>=179 and ll<181) or (cc=172 and ll=180) or (cc=173 and ll=180) or (cc=174 and ll=181) or (cc=175 and ll=181) or (cc=176 and ll>=181 and ll<183) or (cc=177 and ll=182) or (cc=178 and ll=182) or (cc=179 and ll=183) or (cc=180 and ll=183) or (cc=181 and ll=183)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="1000")) then
	if ((cc=118 and ll=162) or (cc=119 and ll>=155 and ll<164) or (cc=120 and ll>=152 and ll<164) or (cc=121 and ll>=152 and ll<165) or (cc=122 and ll>=153 and ll<164) or (cc=123 and ll>=153 and ll<164) or (cc=124 and ll>=154 and ll<165) or (cc=125 and ll>=155 and ll<165) or (cc=126 and ll>=155 and ll<166) or (cc=127 and ll>=156 and ll<167) or (cc=128 and ll>=156 and ll<167) or (cc=129 and ll>=158 and ll<168) or (cc=130 and ll>=159 and ll<168) or (cc=131 and ll>=160 and ll<169) or (cc=132 and ll>=160 and ll<170) or (cc=133 and ll>=161 and ll<171) or (cc=134 and ll>=161 and ll<171) or (cc=135 and ll>=162 and ll<172) or (cc=136 and ll>=163 and ll<172) or (cc=137 and ll>=163 and ll<173) or (cc=138 and ll>=164 and ll<174) or (cc=139 and ll>=166 and ll<174) or (cc=140 and ll>=166 and ll<175) or (cc=141 and ll>=167 and ll<176) or (cc=142 and ll>=168 and ll<176) or (cc=143 and ll>=168 and ll<175) or (cc=144 and ll>=169 and ll<175) or (cc=145 and ll>=170 and ll<176) or (cc=146 and ll>=170 and ll<177) or (cc=147 and ll>=171 and ll<177) or (cc=148 and ll>=172 and ll<178) or (cc=149 and ll>=173 and ll<179) or (cc=150 and ll>=174 and ll<179) or (cc=151 and ll>=174 and ll<180) or (cc=152 and ll>=175 and ll<181) or (cc=153 and ll>=176 and ll<181) or (cc=154 and ll>=176 and ll<182) or (cc=155 and ll>=177 and ll<183) or (cc=156 and ll>=178 and ll<183) or (cc=157 and ll>=178 and ll<184) or (cc=158 and ll>=179 and ll<185) or (cc=159 and ll>=180 and ll<185) or (cc=160 and ll>=181 and ll<186) or (cc=161 and ll>=182 and ll<187) or (cc=162 and ll>=183 and ll<187) or (cc=163 and ll>=183 and ll<188) or (cc=164 and ll>=184 and ll<186) or (cc=165 and ll>=184 and ll<187) or (cc=166 and ll>=185 and ll<188) or (cc=167 and ll>=186 and ll<188) or (cc=168 and ll>=186 and ll<189) or (cc=169 and ll>=187 and ll<190) or (cc=170 and ll=189) or (cc=171 and ll>=189 and ll<191) or (cc=172 and ll=190) or (cc=173 and ll=191) or (cc=174 and ll>=191 and ll<193) or (cc=175 and ll=192) or (cc=176 and ll=193) or (cc=177 and ll>=193 and ll<195) or (cc=178 and ll=194) or (cc=179 and ll=195)) then grbp<="101";
	end if;

elsif ((PT4 ="0001" and PT5 ="1001")) then
	if ((cc=118 and ll=161) or (cc=119 and ll>=157 and ll<162) or (cc=120 and ll>=151 and ll<163) or (cc=121 and ll>=151 and ll<164) or (cc=122 and ll>=152 and ll<163) or (cc=123 and ll>=153 and ll<164) or (cc=124 and ll>=153 and ll<165) or (cc=125 and ll>=154 and ll<165) or (cc=126 and ll>=155 and ll<167) or (cc=127 and ll>=156 and ll<167) or (cc=128 and ll>=157 and ll<168) or (cc=129 and ll>=159 and ll<169) or (cc=130 and ll>=160 and ll<170) or (cc=131 and ll>=161 and ll<171) or (cc=132 and ll>=162 and ll<172) or (cc=133 and ll>=162 and ll<173) or (cc=134 and ll>=163 and ll<174) or (cc=135 and ll>=164 and ll<174) or (cc=136 and ll>=165 and ll<175) or (cc=137 and ll>=166 and ll<176) or (cc=138 and ll>=167 and ll<177) or (cc=139 and ll>=169 and ll<178) or (cc=140 and ll>=170 and ll<179) or (cc=141 and ll>=171 and ll<180) or (cc=142 and ll>=171 and ll<179) or (cc=143 and ll>=172 and ll<179) or (cc=144 and ll>=173 and ll<180) or (cc=145 and ll>=174 and ll<181) or (cc=146 and ll>=175 and ll<182) or (cc=147 and ll>=176 and ll<183) or (cc=148 and ll>=177 and ll<184) or (cc=149 and ll>=179 and ll<185) or (cc=150 and ll>=180 and ll<185) or (cc=151 and ll>=180 and ll<186) or (cc=152 and ll>=182 and ll<187) or (cc=153 and ll>=182 and ll<188) or (cc=154 and ll>=183 and ll<189) or (cc=155 and ll>=184 and ll<190) or (cc=156 and ll>=185 and ll<191) or (cc=157 and ll>=186 and ll<192) or (cc=158 and ll>=188 and ll<193) or (cc=159 and ll>=189 and ll<194) or (cc=160 and ll>=190 and ll<194) or (cc=161 and ll>=191 and ll<195) or (cc=162 and ll>=191 and ll<196) or (cc=163 and ll>=192 and ll<195) or (cc=164 and ll>=193 and ll<196) or (cc=165 and ll>=194 and ll<197) or (cc=166 and ll>=195 and ll<197) or (cc=167 and ll>=196 and ll<198) or (cc=168 and ll=198) or (cc=169 and ll=199) or (cc=170 and ll=200) or (cc=171 and ll>=200 and ll<202) or (cc=172 and ll>=201 and ll<203) or (cc=173 and ll>=202 and ll<204) or (cc=174 and ll>=203 and ll<205) or (cc=175 and ll=204) or (cc=176 and ll=205) or (cc=177 and ll=206)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0000")) then
	if ((cc=118 and ll=159) or (cc=119 and ll>=156 and ll<161) or (cc=120 and ll>=152 and ll<163) or (cc=121 and ll>=150 and ll<161) or (cc=122 and ll>=151 and ll<162) or (cc=123 and ll>=152 and ll<163) or (cc=124 and ll>=153 and ll<165) or (cc=125 and ll>=154 and ll<166) or (cc=126 and ll>=155 and ll<167) or (cc=127 and ll>=156 and ll<168) or (cc=128 and ll>=157 and ll<169) or (cc=129 and ll>=160 and ll<170) or (cc=130 and ll>=161 and ll<171) or (cc=131 and ll>=162 and ll<173) or (cc=132 and ll>=163 and ll<174) or (cc=133 and ll>=164 and ll<175) or (cc=134 and ll>=165 and ll<176) or (cc=135 and ll>=166 and ll<177) or (cc=136 and ll>=167 and ll<178) or (cc=137 and ll>=169 and ll<180) or (cc=138 and ll>=171 and ll<181) or (cc=139 and ll>=172 and ll<182) or (cc=140 and ll>=173 and ll<183) or (cc=141 and ll>=175 and ll<182) or (cc=142 and ll>=176 and ll<183) or (cc=143 and ll>=177 and ll<184) or (cc=144 and ll>=178 and ll<186) or (cc=145 and ll>=179 and ll<187) or (cc=146 and ll>=180 and ll<188) or (cc=147 and ll>=181 and ll<189) or (cc=148 and ll>=184 and ll<190) or (cc=149 and ll>=185 and ll<191) or (cc=150 and ll>=186 and ll<192) or (cc=151 and ll>=187 and ll<194) or (cc=152 and ll>=188 and ll<195) or (cc=153 and ll>=190 and ll<196) or (cc=154 and ll>=191 and ll<197) or (cc=155 and ll>=192 and ll<198) or (cc=156 and ll>=193 and ll<199) or (cc=157 and ll>=195 and ll<201) or (cc=158 and ll>=196 and ll<202) or (cc=159 and ll>=197 and ll<203) or (cc=160 and ll>=198 and ll<203) or (cc=161 and ll>=200 and ll<203) or (cc=162 and ll>=201 and ll<204) or (cc=163 and ll>=202 and ll<205) or (cc=164 and ll>=203 and ll<206) or (cc=165 and ll>=204 and ll<207) or (cc=166 and ll=207) or (cc=167 and ll=208) or (cc=168 and ll>=209 and ll<211) or (cc=169 and ll>=210 and ll<212) or (cc=170 and ll>=211 and ll<213) or (cc=171 and ll>=212 and ll<214) or (cc=172 and ll=214) or (cc=173 and ll=215) or (cc=174 and ll>=216 and ll<218)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0001")) then
	if ((cc=118 and ll=158) or (cc=119 and ll>=156 and ll<160) or (cc=120 and ll>=152 and ll<162) or (cc=121 and ll>=150 and ll<161) or (cc=122 and ll>=149 and ll<162) or (cc=123 and ll>=151 and ll<164) or (cc=124 and ll>=152 and ll<165) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=155 and ll<168) or (cc=127 and ll>=157 and ll<170) or (cc=128 and ll>=158 and ll<171) or (cc=129 and ll>=160 and ll<172) or (cc=130 and ll>=162 and ll<174) or (cc=131 and ll>=163 and ll<175) or (cc=132 and ll>=165 and ll<177) or (cc=133 and ll>=166 and ll<178) or (cc=134 and ll>=168 and ll<179) or (cc=135 and ll>=169 and ll<181) or (cc=136 and ll>=171 and ll<182) or (cc=137 and ll>=172 and ll<184) or (cc=138 and ll>=175 and ll<185) or (cc=139 and ll>=176 and ll<186) or (cc=140 and ll>=177 and ll<185) or (cc=141 and ll>=179 and ll<187) or (cc=142 and ll>=180 and ll<188) or (cc=143 and ll>=182 and ll<190) or (cc=144 and ll>=183 and ll<191) or (cc=145 and ll>=185 and ll<193) or (cc=146 and ll>=188 and ll<194) or (cc=147 and ll>=189 and ll<195) or (cc=148 and ll>=191 and ll<197) or (cc=149 and ll>=192 and ll<198) or (cc=150 and ll>=194 and ll<200) or (cc=151 and ll>=195 and ll<201) or (cc=152 and ll>=196 and ll<203) or (cc=153 and ll>=198 and ll<204) or (cc=154 and ll>=199 and ll<206) or (cc=155 and ll>=202 and ll<207) or (cc=156 and ll>=203 and ll<209) or (cc=157 and ll>=204 and ll<210) or (cc=158 and ll>=206 and ll<209) or (cc=159 and ll>=207 and ll<211) or (cc=160 and ll>=209 and ll<212) or (cc=161 and ll>=210 and ll<214) or (cc=162 and ll>=212 and ll<215) or (cc=163 and ll>=213 and ll<216) or (cc=164 and ll>=216 and ll<218) or (cc=165 and ll>=217 and ll<219) or (cc=166 and ll>=219 and ll<221) or (cc=167 and ll>=220 and ll<222) or (cc=168 and ll>=221 and ll<224) or (cc=169 and ll>=223 and ll<225) or (cc=170 and ll>=224 and ll<227) or (cc=171 and ll>=226 and ll<228)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0010")) then
	if ((cc=119 and ll>=155 and ll<159) or (cc=120 and ll>=153 and ll<161) or (cc=121 and ll>=151 and ll<160) or (cc=122 and ll>=148 and ll<161) or (cc=123 and ll>=149 and ll<163) or (cc=124 and ll>=151 and ll<165) or (cc=125 and ll>=153 and ll<167) or (cc=126 and ll>=154 and ll<169) or (cc=127 and ll>=156 and ll<171) or (cc=128 and ll>=158 and ll<172) or (cc=129 and ll>=161 and ll<174) or (cc=130 and ll>=163 and ll<176) or (cc=131 and ll>=165 and ll<178) or (cc=132 and ll>=166 and ll<179) or (cc=133 and ll>=168 and ll<181) or (cc=134 and ll>=170 and ll<183) or (cc=135 and ll>=172 and ll<185) or (cc=136 and ll>=174 and ll<187) or (cc=137 and ll>=177 and ll<189) or (cc=138 and ll>=178 and ll<188) or (cc=139 and ll>=180 and ll<189) or (cc=140 and ll>=182 and ll<191) or (cc=141 and ll>=184 and ll<193) or (cc=142 and ll>=186 and ll<195) or (cc=143 and ll>=188 and ll<197) or (cc=144 and ll>=189 and ll<199) or (cc=145 and ll>=193 and ll<200) or (cc=146 and ll>=195 and ll<202) or (cc=147 and ll>=196 and ll<204) or (cc=148 and ll>=198 and ll<205) or (cc=149 and ll>=200 and ll<207) or (cc=150 and ll>=201 and ll<209) or (cc=151 and ll>=203 and ll<211) or (cc=152 and ll>=205 and ll<213) or (cc=153 and ll>=208 and ll<215) or (cc=154 and ll>=210 and ll<216) or (cc=155 and ll>=212 and ll<217) or (cc=156 and ll>=213 and ll<217) or (cc=157 and ll>=215 and ll<219) or (cc=158 and ll>=217 and ll<220) or (cc=159 and ll>=219 and ll<222) or (cc=160 and ll>=221 and ll<224) or (cc=161 and ll>=224 and ll<226) or (cc=162 and ll>=225 and ll<228) or (cc=163 and ll>=227 and ll<230) or (cc=164 and ll>=229 and ll<232) or (cc=165 and ll>=231 and ll<233) or (cc=166 and ll>=233 and ll<235) or (cc=167 and ll>=235 and ll<237)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0011")) then
	if ((cc=119 and ll>=154 and ll<158) or (cc=120 and ll>=152 and ll<160) or (cc=121 and ll>=150 and ll<158) or (cc=122 and ll>=148 and ll<161) or (cc=123 and ll>=148 and ll<163) or (cc=124 and ll>=150 and ll<165) or (cc=125 and ll>=151 and ll<167) or (cc=126 and ll>=154 and ll<170) or (cc=127 and ll>=156 and ll<172) or (cc=128 and ll>=158 and ll<174) or (cc=129 and ll>=163 and ll<176) or (cc=130 and ll>=164 and ll<179) or (cc=131 and ll>=166 and ll<181) or (cc=132 and ll>=168 and ll<183) or (cc=133 and ll>=171 and ll<185) or (cc=134 and ll>=173 and ll<187) or (cc=135 and ll>=175 and ll<190) or (cc=136 and ll>=179 and ll<191) or (cc=137 and ll>=181 and ll<191) or (cc=138 and ll>=183 and ll<193) or (cc=139 and ll>=185 and ll<196) or (cc=140 and ll>=188 and ll<198) or (cc=141 and ll>=190 and ll<200) or (cc=142 and ll>=192 and ll<202) or (cc=143 and ll>=196 and ll<205) or (cc=144 and ll>=198 and ll<207) or (cc=145 and ll>=200 and ll<209) or (cc=146 and ll>=202 and ll<211) or (cc=147 and ll>=205 and ll<213) or (cc=148 and ll>=207 and ll<216) or (cc=149 and ll>=209 and ll<218) or (cc=150 and ll>=213 and ll<220) or (cc=151 and ll>=215 and ll<222) or (cc=152 and ll>=217 and ll<221) or (cc=153 and ll>=219 and ll<223) or (cc=154 and ll>=222 and ll<225) or (cc=155 and ll>=224 and ll<228) or (cc=156 and ll>=226 and ll<230) or (cc=157 and ll>=230 and ll<232) or (cc=158 and ll>=232 and ll<234) or (cc=159 and ll>=234 and ll<237) or (cc=160 and ll>=236 and ll<239) or (cc=161 and ll>=239 and ll<241) or (cc=162 and ll>=241 and ll<243) or (cc=163 and ll>=243 and ll<246)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0100")) then
	if ((cc=119 and ll>=154 and ll<156) or (cc=120 and ll>=153 and ll<158) or (cc=121 and ll>=150 and ll<159) or (cc=122 and ll>=149 and ll<160) or (cc=123 and ll>=147 and ll<163) or (cc=124 and ll>=148 and ll<166) or (cc=125 and ll>=151 and ll<169) or (cc=126 and ll>=153 and ll<171) or (cc=127 and ll>=156 and ll<174) or (cc=128 and ll>=159 and ll<177) or (cc=129 and ll>=163 and ll<180) or (cc=130 and ll>=166 and ll<183) or (cc=131 and ll>=169 and ll<185) or (cc=132 and ll>=171 and ll<188) or (cc=133 and ll>=174 and ll<191) or (cc=134 and ll>=177 and ll<193) or (cc=135 and ll>=182 and ll<193) or (cc=136 and ll>=184 and ll<195) or (cc=137 and ll>=186 and ll<199) or (cc=138 and ll>=190 and ll<201) or (cc=139 and ll>=192 and ll<203) or (cc=140 and ll>=195 and ll<207) or (cc=141 and ll>=199 and ll<209) or (cc=142 and ll>=202 and ll<212) or (cc=143 and ll>=205 and ll<215) or (cc=144 and ll>=207 and ll<217) or (cc=145 and ll>=210 and ll<220) or (cc=146 and ll>=213 and ll<223) or (cc=147 and ll>=218 and ll<225) or (cc=148 and ll>=220 and ll<228) or (cc=149 and ll>=223 and ll<228) or (cc=150 and ll>=226 and ll<230) or (cc=151 and ll>=229 and ll<233) or (cc=152 and ll>=231 and ll<236) or (cc=153 and ll>=234 and ll<239) or (cc=154 and ll>=238 and ll<241) or (cc=155 and ll>=241 and ll<244) or (cc=156 and ll>=244 and ll<247) or (cc=157 and ll>=246 and ll<250) or (cc=158 and ll>=250 and ll<252) or (cc=159 and ll=252)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0101")) then
	if ((cc=119 and ll=153) or (cc=120 and ll>=152 and ll<157) or (cc=121 and ll>=151 and ll<158) or (cc=122 and ll>=149 and ll<160) or (cc=123 and ll>=148 and ll<163) or (cc=124 and ll>=147 and ll<166) or (cc=125 and ll>=149 and ll<170) or (cc=126 and ll>=152 and ll<173) or (cc=127 and ll>=156 and ll<177) or (cc=128 and ll>=159 and ll<180) or (cc=129 and ll>=165 and ll<184) or (cc=130 and ll>=168 and ll<187) or (cc=131 and ll>=172 and ll<191) or (cc=132 and ll>=174 and ll<194) or (cc=133 and ll>=178 and ll<195) or (cc=134 and ll>=184 and ll<197) or (cc=135 and ll>=187 and ll<201) or (cc=136 and ll>=190 and ll<204) or (cc=137 and ll>=194 and ll<208) or (cc=138 and ll>=197 and ll<211) or (cc=139 and ll>=203 and ll<215) or (cc=140 and ll>=207 and ll<218) or (cc=141 and ll>=210 and ll<222) or (cc=142 and ll>=213 and ll<225) or (cc=143 and ll>=217 and ll<229) or (cc=144 and ll>=222 and ll<232) or (cc=145 and ll>=225 and ll<231) or (cc=146 and ll>=229 and ll<234) or (cc=147 and ll>=232 and ll<238) or (cc=148 and ll>=236 and ll<241) or (cc=149 and ll>=239 and ll<245) or (cc=150 and ll>=245 and ll<248) or (cc=151 and ll>=248 and ll<252) or (cc=152 and ll>=252 and ll<255) or (cc=153 and ll>=255 and ll<259) or (cc=154 and ll=259)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0110")) then
	if ((cc=120 and ll>=152 and ll<155) or (cc=121 and ll>=151 and ll<157) or (cc=122 and ll>=150 and ll<159) or (cc=123 and ll>=148 and ll<164) or (cc=124 and ll>=147 and ll<168) or (cc=125 and ll>=147 and ll<173) or (cc=126 and ll>=151 and ll<177) or (cc=127 and ll>=155 and ll<182) or (cc=128 and ll>=160 and ll<186) or (cc=129 and ll>=167 and ll<190) or (cc=130 and ll>=171 and ll<195) or (cc=131 and ll>=175 and ll<196) or (cc=132 and ll>=179 and ll<199) or (cc=133 and ll>=186 and ll<203) or (cc=134 and ll>=191 and ll<207) or (cc=135 and ll>=195 and ll<212) or (cc=136 and ll>=200 and ll<217) or (cc=137 and ll>=207 and ll<221) or (cc=138 and ll>=211 and ll<226) or (cc=139 and ll>=216 and ll<230) or (cc=140 and ll>=220 and ll<235) or (cc=141 and ll>=227 and ll<236) or (cc=142 and ll>=232 and ll<239) or (cc=143 and ll>=236 and ll<243) or (cc=144 and ll>=241 and ll<248) or (cc=145 and ll>=248 and ll<252) or (cc=146 and ll>=252 and ll<257) or (cc=147 and ll>=257 and ll<260) or (cc=148 and ll>=260 and ll<265)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="0111")) then
	if ((cc=120 and ll>=150 and ll<152) or (cc=121 and ll>=150 and ll<156) or (cc=122 and ll>=149 and ll<158) or (cc=123 and ll>=149 and ll<164) or (cc=124 and ll>=148 and ll<170) or (cc=125 and ll>=147 and ll<176) or (cc=126 and ll>=147 and ll<182) or (cc=127 and ll>=154 and ll<189) or (cc=128 and ll>=159 and ll<195) or (cc=129 and ll>=169 and ll<197) or (cc=130 and ll>=175 and ll<201) or (cc=131 and ll>=182 and ll<206) or (cc=132 and ll>=190 and ll<213) or (cc=133 and ll>=196 and ll<219) or (cc=134 and ll>=203 and ll<225) or (cc=135 and ll>=212 and ll<231) or (cc=136 and ll>=218 and ll<237) or (cc=137 and ll>=224 and ll<239) or (cc=138 and ll>=234 and ll<243) or (cc=139 and ll>=239 and ll<248) or (cc=140 and ll>=245 and ll<255) or (cc=141 and ll>=255 and ll<261) or (cc=142 and ll>=261 and ll<267) or (cc=143 and ll>=267 and ll<269)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="1000")) then
	if ((cc=121 and ll>=150 and ll<155) or (cc=122 and ll>=149 and ll<156) or (cc=123 and ll>=149 and ll<166) or (cc=124 and ll>=148 and ll<175) or (cc=125 and ll>=148 and ll<184) or (cc=126 and ll>=147 and ll<193) or (cc=127 and ll>=151 and ll<198) or (cc=128 and ll>=160 and ll<202) or (cc=129 and ll>=174 and ll<211) or (cc=130 and ll>=184 and ll<221) or (cc=131 and ll>=197 and ll<230) or (cc=132 and ll>=206 and ll<240) or (cc=133 and ll>=220 and ll<241) or (cc=134 and ll>=234 and ll<249) or (cc=135 and ll>=244 and ll<258) or (cc=136 and ll>=258 and ll<268) or (cc=137 and ll>=268 and ll<272)) then grbp<="101";
	end if;

elsif ((PT4 ="0010" and PT5 ="1001")) then
	if ((cc=121 and ll>=149 and ll<152) or (cc=122 and ll>=149 and ll<155) or (cc=123 and ll>=148 and ll<170) or (cc=124 and ll>=148 and ll<188) or (cc=125 and ll>=148 and ll<198) or (cc=126 and ll>=148 and ll<207) or (cc=127 and ll>=148 and ll<225) or (cc=128 and ll>=160 and ll<242) or (cc=129 and ll>=197 and ll<244) or (cc=130 and ll>=225 and ll<262) or (cc=131 and ll>=262 and ll<274)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0000")) then
	if ((cc=122 and ll>=148 and ll<154) or (cc=123 and ll>=148 and ll<198) or (cc=124 and ll>=148 and ll<242) or (cc=125 and ll>=148 and ll<275) or (cc=126 and ll>=148 and ll<253) or (cc=127 and ll>=148 and ll<209) or (cc=128 and ll>=161 and ll<165)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0001")) then
	if ((cc=119 and ll>=268 and ll<274) or (cc=120 and ll>=229 and ll<268) or (cc=121 and ll>=189 and ll<253) or (cc=122 and ll>=150 and ll<239) or (cc=123 and ll>=147 and ll<229) or (cc=124 and ll>=148 and ll<210) or (cc=125 and ll>=148 and ll<200) or (cc=126 and ll>=148 and ll<187) or (cc=127 and ll>=148 and ll<170) or (cc=128 and ll>=148 and ll<161)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0010")) then
	if ((cc=113 and ll>=271 and ll<273) or (cc=114 and ll>=261 and ll<271) or (cc=115 and ll>=251 and ll<261) or (cc=116 and ll>=232 and ll<251) or (cc=117 and ll>=222 and ll<246) or (cc=118 and ll>=212 and ll<238) or (cc=119 and ll>=193 and ll<230) or (cc=120 and ll>=184 and ll<223) or (cc=121 and ll>=175 and ll<213) or (cc=122 and ll>=165 and ll<209) or (cc=123 and ll>=147 and ll<199) or (cc=124 and ll>=147 and ll<190) or (cc=125 and ll>=148 and ll<185) or (cc=126 and ll>=148 and ll<176) or (cc=127 and ll>=148 and ll<166) or (cc=128 and ll>=149 and ll<161) or (cc=129 and ll>=149 and ll<151)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0011")) then
	if ((cc=108 and ll>=263 and ll<270) or (cc=109 and ll>=257 and ll<263) or (cc=110 and ll>=250 and ll<257) or (cc=111 and ll>=245 and ll<250) or (cc=112 and ll>=232 and ll<248) or (cc=113 and ll>=225 and ll<241) or (cc=114 and ll>=219 and ll<236) or (cc=115 and ll>=213 and ll<229) or (cc=116 and ll>=207 and ll<226) or (cc=117 and ll>=194 and ll<220) or (cc=118 and ll>=188 and ll<214) or (cc=119 and ll>=182 and ll<208) or (cc=120 and ll>=175 and ll<205) or (cc=121 and ll>=169 and ll<198) or (cc=122 and ll>=163 and ll<192) or (cc=123 and ll>=151 and ll<187) or (cc=124 and ll>=147 and ll<183) or (cc=125 and ll>=147 and ll<177) or (cc=126 and ll>=148 and ll<171) or (cc=127 and ll>=149 and ll<166) or (cc=128 and ll>=149 and ll<162) or (cc=129 and ll>=150 and ll<155)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0100")) then
	if ((cc=102 and ll>=262 and ll<265) or (cc=103 and ll>=258 and ll<263) or (cc=104 and ll>=253 and ll<258) or (cc=105 and ll>=249 and ll<253) or (cc=106 and ll>=244 and ll<249) or (cc=107 and ll>=240 and ll<246) or (cc=108 and ll>=231 and ll<242) or (cc=109 and ll>=226 and ll<238) or (cc=110 and ll>=221 and ll<234) or (cc=111 and ll>=217 and ll<229) or (cc=112 and ll>=212 and ll<226) or (cc=113 and ll>=208 and ll<222) or (cc=114 and ll>=203 and ll<218) or (cc=115 and ll>=199 and ll<213) or (cc=116 and ll>=189 and ll<208) or (cc=117 and ll>=185 and ll<206) or (cc=118 and ll>=180 and ll<202) or (cc=119 and ll>=176 and ll<198) or (cc=120 and ll>=171 and ll<193) or (cc=121 and ll>=167 and ll<189) or (cc=122 and ll>=162 and ll<186) or (cc=123 and ll>=157 and ll<182) or (cc=124 and ll>=148 and ll<177) or (cc=125 and ll>=147 and ll<173) or (cc=126 and ll>=147 and ll<168) or (cc=127 and ll>=148 and ll<166) or (cc=128 and ll>=149 and ll<161) or (cc=129 and ll>=150 and ll<157) or (cc=130 and ll>=151 and ll<153)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0101")) then
	if ((cc=97 and ll>=256 and ll<260) or (cc=98 and ll>=253 and ll<256) or (cc=99 and ll>=249 and ll<253) or (cc=100 and ll>=246 and ll<250) or (cc=101 and ll>=242 and ll<246) or (cc=102 and ll>=239 and ll<243) or (cc=103 and ll>=235 and ll<241) or (cc=104 and ll>=228 and ll<238) or (cc=105 and ll>=224 and ll<234) or (cc=106 and ll>=221 and ll<231) or (cc=107 and ll>=217 and ll<227) or (cc=108 and ll>=214 and ll<224) or (cc=109 and ll>=210 and ll<222) or (cc=110 and ll>=207 and ll<218) or (cc=111 and ll>=203 and ll<215) or (cc=112 and ll>=200 and ll<211) or (cc=113 and ll>=196 and ll<208) or (cc=114 and ll>=189 and ll<205) or (cc=115 and ll>=186 and ll<203) or (cc=116 and ll>=182 and ll<200) or (cc=117 and ll>=179 and ll<196) or (cc=118 and ll>=175 and ll<193) or (cc=119 and ll>=172 and ll<189) or (cc=120 and ll>=168 and ll<186) or (cc=121 and ll>=165 and ll<185) or (cc=122 and ll>=161 and ll<181) or (cc=123 and ll>=158 and ll<178) or (cc=124 and ll>=150 and ll<174) or (cc=125 and ll>=147 and ll<170) or (cc=126 and ll>=148 and ll<167) or (cc=127 and ll>=149 and ll<165) or (cc=128 and ll>=150 and ll<162) or (cc=129 and ll>=151 and ll<158) or (cc=130 and ll>=152 and ll<155)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0110")) then
	if ((cc=92 and ll>=251 and ll<253) or (cc=93 and ll>=248 and ll<251) or (cc=94 and ll>=245 and ll<248) or (cc=95 and ll>=242 and ll<245) or (cc=96 and ll>=239 and ll<242) or (cc=97 and ll>=237 and ll<240) or (cc=98 and ll>=234 and ll<237) or (cc=99 and ll>=231 and ll<235) or (cc=100 and ll>=225 and ll<233) or (cc=101 and ll>=222 and ll<231) or (cc=102 and ll>=220 and ll<227) or (cc=103 and ll>=216 and ll<225) or (cc=104 and ll>=214 and ll<222) or (cc=105 and ll>=211 and ll<219) or (cc=106 and ll>=208 and ll<218) or (cc=107 and ll>=206 and ll<216) or (cc=108 and ll>=203 and ll<212) or (cc=109 and ll>=200 and ll<210) or (cc=110 and ll>=197 and ll<207) or (cc=111 and ll>=195 and ll<204) or (cc=112 and ll>=191 and ll<202) or (cc=113 and ll>=185 and ll<200) or (cc=114 and ll>=183 and ll<198) or (cc=115 and ll>=180 and ll<195) or (cc=116 and ll>=177 and ll<192) or (cc=117 and ll>=175 and ll<190) or (cc=118 and ll>=171 and ll<186) or (cc=119 and ll>=169 and ll<184) or (cc=120 and ll>=166 and ll<183) or (cc=121 and ll>=163 and ll<180) or (cc=122 and ll>=161 and ll<177) or (cc=123 and ll>=158 and ll<175) or (cc=124 and ll>=155 and ll<171) or (cc=125 and ll>=148 and ll<169) or (cc=126 and ll>=147 and ll<167) or (cc=127 and ll>=148 and ll<165) or (cc=128 and ll>=149 and ll<162) or (cc=129 and ll>=150 and ll<159) or (cc=130 and ll>=152 and ll<157) or (cc=131 and ll=153)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="0111")) then
	if ((cc=87 and ll>=244 and ll<246) or (cc=88 and ll>=242 and ll<244) or (cc=89 and ll>=240 and ll<242) or (cc=90 and ll>=238 and ll<240) or (cc=91 and ll>=235 and ll<238) or (cc=92 and ll>=233 and ll<236) or (cc=93 and ll>=231 and ll<233) or (cc=94 and ll>=229 and ll<231) or (cc=95 and ll>=226 and ll<230) or (cc=96 and ll>=224 and ll<228) or (cc=97 and ll>=219 and ll<226) or (cc=98 and ll>=217 and ll<224) or (cc=99 and ll>=215 and ll<221) or (cc=100 and ll>=212 and ll<219) or (cc=101 and ll>=210 and ll<217) or (cc=102 and ll>=208 and ll<215) or (cc=103 and ll>=206 and ll<214) or (cc=104 and ll>=203 and ll<212) or (cc=105 and ll>=201 and ll<209) or (cc=106 and ll>=199 and ll<207) or (cc=107 and ll>=197 and ll<205) or (cc=108 and ll>=194 and ll<203) or (cc=109 and ll>=192 and ll<200) or (cc=110 and ll>=190 and ll<199) or (cc=111 and ll>=185 and ll<197) or (cc=112 and ll>=183 and ll<195) or (cc=113 and ll>=180 and ll<193) or (cc=114 and ll>=178 and ll<191) or (cc=115 and ll>=176 and ll<188) or (cc=116 and ll>=174 and ll<186) or (cc=117 and ll>=171 and ll<184) or (cc=118 and ll>=169 and ll<183) or (cc=119 and ll>=167 and ll<181) or (cc=120 and ll>=165 and ll<179) or (cc=121 and ll>=163 and ll<176) or (cc=122 and ll>=160 and ll<174) or (cc=123 and ll>=158 and ll<172) or (cc=124 and ll>=156 and ll<170) or (cc=125 and ll>=150 and ll<167) or (cc=126 and ll>=148 and ll<167) or (cc=127 and ll>=147 and ll<165) or (cc=128 and ll>=148 and ll<163) or (cc=129 and ll>=151 and ll<161) or (cc=130 and ll>=152 and ll<158) or (cc=131 and ll>=154 and ll<156)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="1000")) then
	if ((cc=83 and ll>=236 and ll<238) or (cc=84 and ll>=234 and ll<236) or (cc=85 and ll>=232 and ll<234) or (cc=86 and ll>=230 and ll<232) or (cc=87 and ll=229) or (cc=88 and ll>=227 and ll<229) or (cc=89 and ll>=224 and ll<227) or (cc=90 and ll>=223 and ll<225) or (cc=91 and ll>=221 and ll<224) or (cc=92 and ll>=219 and ll<223) or (cc=93 and ll>=218 and ll<221) or (cc=94 and ll>=213 and ll<219) or (cc=95 and ll>=211 and ll<218) or (cc=96 and ll>=210 and ll<215) or (cc=97 and ll>=208 and ll<213) or (cc=98 and ll>=206 and ll<212) or (cc=99 and ll>=204 and ll<210) or (cc=100 and ll>=202 and ll<210) or (cc=101 and ll>=200 and ll<207) or (cc=102 and ll>=198 and ll<206) or (cc=103 and ll>=197 and ll<204) or (cc=104 and ll>=195 and ll<202) or (cc=105 and ll>=193 and ll<201) or (cc=106 and ll>=191 and ll<199) or (cc=107 and ll>=189 and ll<197) or (cc=108 and ll>=187 and ll<195) or (cc=109 and ll>=186 and ll<195) or (cc=110 and ll>=181 and ll<193) or (cc=111 and ll>=179 and ll<191) or (cc=112 and ll>=178 and ll<189) or (cc=113 and ll>=176 and ll<187) or (cc=114 and ll>=174 and ll<185) or (cc=115 and ll>=172 and ll<184) or (cc=116 and ll>=170 and ll<182) or (cc=117 and ll>=168 and ll<181) or (cc=118 and ll>=166 and ll<179) or (cc=119 and ll>=165 and ll<178) or (cc=120 and ll>=163 and ll<176) or (cc=121 and ll>=161 and ll<174) or (cc=122 and ll>=160 and ll<173) or (cc=123 and ll>=158 and ll<171) or (cc=124 and ll>=156 and ll<169) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=150 and ll<167) or (cc=127 and ll>=147 and ll<165) or (cc=128 and ll>=149 and ll<163) or (cc=129 and ll>=150 and ll<161) or (cc=130 and ll>=153 and ll<159) or (cc=131 and ll>=155 and ll<157)) then grbp<="101";
	end if;

elsif ((PT4 ="0011" and PT5 ="1001")) then
	if ((cc=79 and ll=227) or (cc=80 and ll=226) or (cc=81 and ll>=224 and ll<226) or (cc=82 and ll=223) or (cc=83 and ll>=221 and ll<223) or (cc=84 and ll=220) or (cc=85 and ll>=218 and ll<220) or (cc=86 and ll=217) or (cc=87 and ll>=215 and ll<217) or (cc=88 and ll>=214 and ll<216) or (cc=89 and ll>=212 and ll<216) or (cc=90 and ll>=211 and ll<214) or (cc=91 and ll>=210 and ll<213) or (cc=92 and ll>=206 and ll<211) or (cc=93 and ll>=204 and ll<210) or (cc=94 and ll>=203 and ll<208) or (cc=95 and ll>=201 and ll<207) or (cc=96 and ll>=200 and ll<205) or (cc=97 and ll>=198 and ll<204) or (cc=98 and ll>=197 and ll<203) or (cc=99 and ll>=195 and ll<202) or (cc=100 and ll>=194 and ll<200) or (cc=101 and ll>=192 and ll<199) or (cc=102 and ll>=191 and ll<197) or (cc=103 and ll>=189 and ll<196) or (cc=104 and ll>=188 and ll<195) or (cc=105 and ll>=186 and ll<193) or (cc=106 and ll>=185 and ll<192) or (cc=107 and ll>=183 and ll<192) or (cc=108 and ll>=182 and ll<190) or (cc=109 and ll>=178 and ll<189) or (cc=110 and ll>=177 and ll<187) or (cc=111 and ll>=175 and ll<186) or (cc=112 and ll>=174 and ll<184) or (cc=113 and ll>=172 and ll<183) or (cc=114 and ll>=171 and ll<181) or (cc=115 and ll>=169 and ll<180) or (cc=116 and ll>=168 and ll<180) or (cc=117 and ll>=166 and ll<178) or (cc=118 and ll>=165 and ll<177) or (cc=119 and ll>=163 and ll<175) or (cc=120 and ll>=162 and ll<174) or (cc=121 and ll>=160 and ll<172) or (cc=122 and ll>=159 and ll<171) or (cc=123 and ll>=157 and ll<170) or (cc=124 and ll>=156 and ll<168) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=150 and ll<166) or (cc=127 and ll>=149 and ll<164) or (cc=128 and ll>=148 and ll<163) or (cc=129 and ll>=150 and ll<161) or (cc=130 and ll>=153 and ll<160) or (cc=131 and ll>=155 and ll<159)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0000")) then
	if ((cc=76 and ll=217) or (cc=77 and ll>=215 and ll<217) or (cc=78 and ll>=214 and ll<216) or (cc=79 and ll>=213 and ll<215) or (cc=80 and ll>=212 and ll<214) or (cc=81 and ll=211) or (cc=82 and ll=210) or (cc=83 and ll=209) or (cc=84 and ll>=207 and ll<209) or (cc=85 and ll>=206 and ll<208) or (cc=86 and ll>=205 and ll<208) or (cc=87 and ll>=204 and ll<207) or (cc=88 and ll>=203 and ll<206) or (cc=89 and ll>=199 and ll<205) or (cc=90 and ll>=198 and ll<203) or (cc=91 and ll>=197 and ll<202) or (cc=92 and ll>=196 and ll<201) or (cc=93 and ll>=195 and ll<200) or (cc=94 and ll>=193 and ll<199) or (cc=95 and ll>=192 and ll<198) or (cc=96 and ll>=191 and ll<197) or (cc=97 and ll>=190 and ll<196) or (cc=98 and ll>=189 and ll<195) or (cc=99 and ll>=187 and ll<194) or (cc=100 and ll>=186 and ll<193) or (cc=101 and ll>=185 and ll<191) or (cc=102 and ll>=184 and ll<190) or (cc=103 and ll>=183 and ll<189) or (cc=104 and ll>=182 and ll<188) or (cc=105 and ll>=180 and ll<188) or (cc=106 and ll>=179 and ll<187) or (cc=107 and ll>=178 and ll<186) or (cc=108 and ll>=175 and ll<185) or (cc=109 and ll>=174 and ll<183) or (cc=110 and ll>=173 and ll<182) or (cc=111 and ll>=171 and ll<181) or (cc=112 and ll>=170 and ll<180) or (cc=113 and ll>=169 and ll<179) or (cc=114 and ll>=168 and ll<178) or (cc=115 and ll>=167 and ll<178) or (cc=116 and ll>=166 and ll<177) or (cc=117 and ll>=165 and ll<176) or (cc=118 and ll>=163 and ll<174) or (cc=119 and ll>=162 and ll<173) or (cc=120 and ll>=161 and ll<172) or (cc=121 and ll>=160 and ll<170) or (cc=122 and ll>=159 and ll<169) or (cc=123 and ll>=158 and ll<168) or (cc=124 and ll>=156 and ll<167) or (cc=125 and ll>=155 and ll<167) or (cc=126 and ll>=154 and ll<166) or (cc=127 and ll>=150 and ll<165) or (cc=128 and ll>=149 and ll<164) or (cc=129 and ll>=149 and ll<162) or (cc=130 and ll>=152 and ll<161) or (cc=131 and ll>=156 and ll<160)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0001")) then
	if ((cc=73 and ll>=206 and ll<208) or (cc=74 and ll=206) or (cc=75 and ll=205) or (cc=76 and ll=204) or (cc=77 and ll=203) or (cc=78 and ll>=202 and ll<204) or (cc=79 and ll=201) or (cc=80 and ll>=200 and ll<202) or (cc=81 and ll>=199 and ll<201) or (cc=82 and ll=199) or (cc=83 and ll>=198 and ll<200) or (cc=84 and ll>=197 and ll<199) or (cc=85 and ll>=196 and ll<198) or (cc=86 and ll>=195 and ll<198) or (cc=87 and ll>=194 and ll<196) or (cc=88 and ll>=191 and ll<196) or (cc=89 and ll>=190 and ll<195) or (cc=90 and ll>=189 and ll<194) or (cc=91 and ll>=188 and ll<193) or (cc=92 and ll>=187 and ll<192) or (cc=93 and ll>=186 and ll<192) or (cc=94 and ll>=185 and ll<191) or (cc=95 and ll>=184 and ll<190) or (cc=96 and ll>=184 and ll<189) or (cc=97 and ll>=183 and ll<189) or (cc=98 and ll>=182 and ll<188) or (cc=99 and ll>=181 and ll<187) or (cc=100 and ll>=180 and ll<186) or (cc=101 and ll>=179 and ll<185) or (cc=102 and ll>=178 and ll<184) or (cc=103 and ll>=177 and ll<183) or (cc=104 and ll>=177 and ll<183) or (cc=105 and ll>=175 and ll<183) or (cc=106 and ll>=175 and ll<182) or (cc=107 and ll>=172 and ll<181) or (cc=108 and ll>=171 and ll<180) or (cc=109 and ll>=170 and ll<179) or (cc=110 and ll>=169 and ll<178) or (cc=111 and ll>=168 and ll<177) or (cc=112 and ll>=167 and ll<176) or (cc=113 and ll>=166 and ll<175) or (cc=114 and ll>=165 and ll<175) or (cc=115 and ll>=165 and ll<174) or (cc=116 and ll>=163 and ll<174) or (cc=117 and ll>=163 and ll<173) or (cc=118 and ll>=162 and ll<172) or (cc=119 and ll>=161 and ll<171) or (cc=120 and ll>=160 and ll<170) or (cc=121 and ll>=159 and ll<169) or (cc=122 and ll>=158 and ll<168) or (cc=123 and ll>=157 and ll<168) or (cc=124 and ll>=156 and ll<167) or (cc=125 and ll>=156 and ll<167) or (cc=126 and ll>=154 and ll<166) or (cc=127 and ll>=151 and ll<165) or (cc=128 and ll>=150 and ll<164) or (cc=129 and ll>=150 and ll<163) or (cc=130 and ll>=151 and ll<162) or (cc=131 and ll>=156 and ll<161)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0010")) then
	if ((cc=71 and ll>=195 and ll<197) or (cc=72 and ll=195) or (cc=73 and ll=194) or (cc=74 and ll>=193 and ll<195) or (cc=75 and ll=193) or (cc=76 and ll>=192 and ll<194) or (cc=77 and ll=192) or (cc=78 and ll=191) or (cc=79 and ll=190) or (cc=80 and ll>=189 and ll<191) or (cc=81 and ll>=189 and ll<191) or (cc=82 and ll>=188 and ll<190) or (cc=83 and ll>=188 and ll<190) or (cc=84 and ll>=187 and ll<189) or (cc=85 and ll>=186 and ll<189) or (cc=86 and ll>=183 and ll<188) or (cc=87 and ll>=183 and ll<187) or (cc=88 and ll>=182 and ll<187) or (cc=89 and ll>=182 and ll<186) or (cc=90 and ll>=181 and ll<185) or (cc=91 and ll>=180 and ll<184) or (cc=92 and ll>=179 and ll<185) or (cc=93 and ll>=179 and ll<184) or (cc=94 and ll>=178 and ll<184) or (cc=95 and ll>=177 and ll<183) or (cc=96 and ll>=177 and ll<182) or (cc=97 and ll>=176 and ll<182) or (cc=98 and ll>=176 and ll<181) or (cc=99 and ll>=175 and ll<180) or (cc=100 and ll>=174 and ll<180) or (cc=101 and ll>=173 and ll<179) or (cc=102 and ll>=173 and ll<179) or (cc=103 and ll>=172 and ll<179) or (cc=104 and ll>=172 and ll<178) or (cc=105 and ll>=171 and ll<178) or (cc=106 and ll>=170 and ll<177) or (cc=107 and ll>=167 and ll<176) or (cc=108 and ll>=167 and ll<175) or (cc=109 and ll>=166 and ll<175) or (cc=110 and ll>=166 and ll<174) or (cc=111 and ll>=165 and ll<174) or (cc=112 and ll>=164 and ll<173) or (cc=113 and ll>=163 and ll<173) or (cc=114 and ll>=163 and ll<173) or (cc=115 and ll>=162 and ll<172) or (cc=116 and ll>=162 and ll<171) or (cc=117 and ll>=161 and ll<171) or (cc=118 and ll>=160 and ll<170) or (cc=119 and ll>=160 and ll<169) or (cc=120 and ll>=159 and ll<169) or (cc=121 and ll>=158 and ll<168) or (cc=122 and ll>=157 and ll<167) or (cc=123 and ll>=157 and ll<167) or (cc=124 and ll>=156 and ll<167) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=155 and ll<166) or (cc=127 and ll>=152 and ll<165) or (cc=128 and ll>=151 and ll<164) or (cc=129 and ll>=151 and ll<164) or (cc=130 and ll>=151 and ll<163) or (cc=131 and ll>=156 and ll<163)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0011")) then
	if ((cc=69 and ll=184) or (cc=70 and ll=184) or (cc=71 and ll=183) or (cc=72 and ll=183) or (cc=73 and ll>=182 and ll<184) or (cc=74 and ll=182) or (cc=75 and ll=182) or (cc=76 and ll=181) or (cc=77 and ll=181) or (cc=78 and ll>=180 and ll<182) or (cc=79 and ll=180) or (cc=80 and ll>=179 and ll<181) or (cc=81 and ll>=179 and ll<181) or (cc=82 and ll>=178 and ll<181) or (cc=83 and ll>=178 and ll<180) or (cc=84 and ll>=178 and ll<180) or (cc=85 and ll>=175 and ll<180) or (cc=86 and ll>=175 and ll<179) or (cc=87 and ll>=174 and ll<179) or (cc=88 and ll>=174 and ll<178) or (cc=89 and ll>=173 and ll<178) or (cc=90 and ll>=173 and ll<177) or (cc=91 and ll>=173 and ll<178) or (cc=92 and ll>=172 and ll<177) or (cc=93 and ll>=172 and ll<177) or (cc=94 and ll>=171 and ll<177) or (cc=95 and ll>=171 and ll<176) or (cc=96 and ll>=170 and ll<176) or (cc=97 and ll>=170 and ll<175) or (cc=98 and ll>=169 and ll<175) or (cc=99 and ll>=169 and ll<174) or (cc=100 and ll>=169 and ll<174) or (cc=101 and ll>=168 and ll<174) or (cc=102 and ll>=168 and ll<174) or (cc=103 and ll>=167 and ll<174) or (cc=104 and ll>=167 and ll<173) or (cc=105 and ll>=167 and ll<173) or (cc=106 and ll>=164 and ll<172) or (cc=107 and ll>=164 and ll<172) or (cc=108 and ll>=163 and ll<172) or (cc=109 and ll>=163 and ll<171) or (cc=110 and ll>=162 and ll<171) or (cc=111 and ll>=162 and ll<170) or (cc=112 and ll>=161 and ll<170) or (cc=113 and ll>=161 and ll<170) or (cc=114 and ll>=161 and ll<170) or (cc=115 and ll>=160 and ll<170) or (cc=116 and ll>=160 and ll<169) or (cc=117 and ll>=159 and ll<169) or (cc=118 and ll>=159 and ll<168) or (cc=119 and ll>=158 and ll<168) or (cc=120 and ll>=158 and ll<167) or (cc=121 and ll>=158 and ll<167) or (cc=122 and ll>=157 and ll<167) or (cc=123 and ll>=157 and ll<166) or (cc=124 and ll>=156 and ll<167) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=155 and ll<166) or (cc=127 and ll>=155 and ll<165) or (cc=128 and ll>=152 and ll<165) or (cc=129 and ll>=152 and ll<164) or (cc=130 and ll>=152 and ll<164) or (cc=131 and ll>=156 and ll<164)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0100")) then
	if ((cc=68 and ll=172) or (cc=69 and ll=172) or (cc=70 and ll=172) or (cc=71 and ll=172) or (cc=72 and ll>=171 and ll<173) or (cc=73 and ll=171) or (cc=74 and ll=171) or (cc=75 and ll=171) or (cc=76 and ll=171) or (cc=77 and ll>=170 and ll<172) or (cc=78 and ll=170) or (cc=79 and ll>=170 and ll<172) or (cc=80 and ll>=170 and ll<172) or (cc=81 and ll>=170 and ll<172) or (cc=82 and ll>=169 and ll<171) or (cc=83 and ll>=169 and ll<171) or (cc=84 and ll>=169 and ll<171) or (cc=85 and ll>=167 and ll<171) or (cc=86 and ll>=166 and ll<171) or (cc=87 and ll>=166 and ll<170) or (cc=88 and ll>=166 and ll<170) or (cc=89 and ll>=166 and ll<170) or (cc=90 and ll>=166 and ll<171) or (cc=91 and ll>=165 and ll<170) or (cc=92 and ll>=165 and ll<170) or (cc=93 and ll>=165 and ll<170) or (cc=94 and ll>=165 and ll<170) or (cc=95 and ll>=165 and ll<170) or (cc=96 and ll>=164 and ll<169) or (cc=97 and ll>=164 and ll<169) or (cc=98 and ll>=164 and ll<169) or (cc=99 and ll>=164 and ll<169) or (cc=100 and ll>=163 and ll<169) or (cc=101 and ll>=163 and ll<169) or (cc=102 and ll>=163 and ll<169) or (cc=103 and ll>=163 and ll<169) or (cc=104 and ll>=163 and ll<169) or (cc=105 and ll>=162 and ll<168) or (cc=106 and ll>=160 and ll<168) or (cc=107 and ll>=160 and ll<168) or (cc=108 and ll>=160 and ll<168) or (cc=109 and ll>=159 and ll<168) or (cc=110 and ll>=159 and ll<167) or (cc=111 and ll>=159 and ll<167) or (cc=112 and ll>=159 and ll<168) or (cc=113 and ll>=159 and ll<168) or (cc=114 and ll>=158 and ll<167) or (cc=115 and ll>=158 and ll<167) or (cc=116 and ll>=158 and ll<167) or (cc=117 and ll>=158 and ll<167) or (cc=118 and ll>=157 and ll<167) or (cc=119 and ll>=157 and ll<166) or (cc=120 and ll>=157 and ll<166) or (cc=121 and ll>=157 and ll<166) or (cc=122 and ll>=157 and ll<166) or (cc=123 and ll>=156 and ll<166) or (cc=124 and ll>=156 and ll<166) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=156 and ll<166) or (cc=127 and ll>=155 and ll<166) or (cc=128 and ll>=153 and ll<165) or (cc=129 and ll>=153 and ll<165) or (cc=130 and ll>=153 and ll<165) or (cc=131 and ll>=153 and ll<165)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0101")) then
	if ((cc=68 and ll=160) or (cc=69 and ll=160) or (cc=70 and ll=160) or (cc=71 and ll=160) or (cc=72 and ll=160) or (cc=73 and ll=160) or (cc=74 and ll=160) or (cc=75 and ll=160) or (cc=76 and ll=160) or (cc=77 and ll=160) or (cc=78 and ll=160) or (cc=79 and ll>=160 and ll<162) or (cc=80 and ll>=160 and ll<162) or (cc=81 and ll>=160 and ll<162) or (cc=82 and ll>=160 and ll<162) or (cc=83 and ll>=160 and ll<162) or (cc=84 and ll>=158 and ll<162) or (cc=85 and ll>=158 and ll<162) or (cc=86 and ll>=158 and ll<162) or (cc=87 and ll>=158 and ll<162) or (cc=88 and ll>=158 and ll<162) or (cc=89 and ll>=158 and ll<162) or (cc=90 and ll>=158 and ll<163) or (cc=91 and ll>=158 and ll<163) or (cc=92 and ll>=158 and ll<163) or (cc=93 and ll>=158 and ll<163) or (cc=94 and ll>=158 and ll<163) or (cc=95 and ll>=158 and ll<163) or (cc=96 and ll>=158 and ll<163) or (cc=97 and ll>=158 and ll<163) or (cc=98 and ll>=158 and ll<163) or (cc=99 and ll>=158 and ll<163) or (cc=100 and ll>=158 and ll<163) or (cc=101 and ll>=158 and ll<164) or (cc=102 and ll>=158 and ll<164) or (cc=103 and ll>=158 and ll<164) or (cc=104 and ll>=158 and ll<164) or (cc=105 and ll>=158 and ll<164) or (cc=106 and ll>=156 and ll<164) or (cc=107 and ll>=156 and ll<164) or (cc=108 and ll>=156 and ll<164) or (cc=109 and ll>=156 and ll<164) or (cc=110 and ll>=156 and ll<164) or (cc=111 and ll>=156 and ll<164) or (cc=112 and ll>=156 and ll<165) or (cc=113 and ll>=156 and ll<165) or (cc=114 and ll>=156 and ll<165) or (cc=115 and ll>=156 and ll<165) or (cc=116 and ll>=156 and ll<165) or (cc=117 and ll>=156 and ll<165) or (cc=118 and ll>=156 and ll<165) or (cc=119 and ll>=156 and ll<165) or (cc=120 and ll>=156 and ll<165) or (cc=121 and ll>=156 and ll<165) or (cc=122 and ll>=156 and ll<165) or (cc=123 and ll>=156 and ll<166) or (cc=124 and ll>=156 and ll<166) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=156 and ll<166) or (cc=127 and ll>=156 and ll<166) or (cc=128 and ll>=154 and ll<166) or (cc=129 and ll>=154 and ll<166) or (cc=130 and ll>=154 and ll<166) or (cc=131 and ll>=154 and ll<166)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0110")) then
	if ((cc=68 and ll=149) or (cc=69 and ll=149) or (cc=70 and ll=149) or (cc=71 and ll=149) or (cc=72 and ll=149) or (cc=73 and ll>=149 and ll<151) or (cc=74 and ll=150) or (cc=75 and ll=150) or (cc=76 and ll=150) or (cc=77 and ll=150) or (cc=78 and ll>=150 and ll<152) or (cc=79 and ll>=151 and ll<153) or (cc=80 and ll>=151 and ll<153) or (cc=81 and ll>=151 and ll<153) or (cc=82 and ll>=151 and ll<153) or (cc=83 and ll>=151 and ll<154) or (cc=84 and ll>=152 and ll<154) or (cc=85 and ll>=150 and ll<154) or (cc=86 and ll>=150 and ll<154) or (cc=87 and ll>=150 and ll<154) or (cc=88 and ll>=150 and ll<155) or (cc=89 and ll>=151 and ll<155) or (cc=90 and ll>=151 and ll<156) or (cc=91 and ll>=151 and ll<156) or (cc=92 and ll>=151 and ll<156) or (cc=93 and ll>=151 and ll<157) or (cc=94 and ll>=152 and ll<157) or (cc=95 and ll>=152 and ll<157) or (cc=96 and ll>=152 and ll<157) or (cc=97 and ll>=152 and ll<157) or (cc=98 and ll>=152 and ll<158) or (cc=99 and ll>=153 and ll<158) or (cc=100 and ll>=153 and ll<158) or (cc=101 and ll>=153 and ll<159) or (cc=102 and ll>=153 and ll<159) or (cc=103 and ll>=153 and ll<160) or (cc=104 and ll>=154 and ll<160) or (cc=105 and ll>=154 and ll<160) or (cc=106 and ll>=154 and ll<160) or (cc=107 and ll>=152 and ll<160) or (cc=108 and ll>=153 and ll<161) or (cc=109 and ll>=153 and ll<161) or (cc=110 and ll>=153 and ll<161) or (cc=111 and ll>=153 and ll<161) or (cc=112 and ll>=153 and ll<162) or (cc=113 and ll>=154 and ll<163) or (cc=114 and ll>=154 and ll<163) or (cc=115 and ll>=154 and ll<163) or (cc=116 and ll>=154 and ll<163) or (cc=117 and ll>=154 and ll<163) or (cc=118 and ll>=155 and ll<164) or (cc=119 and ll>=155 and ll<164) or (cc=120 and ll>=155 and ll<164) or (cc=121 and ll>=155 and ll<164) or (cc=122 and ll>=155 and ll<164) or (cc=123 and ll>=156 and ll<166) or (cc=124 and ll>=156 and ll<166) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=156 and ll<166) or (cc=127 and ll>=156 and ll<166) or (cc=128 and ll>=157 and ll<167) or (cc=129 and ll>=155 and ll<167) or (cc=130 and ll>=155 and ll<167) or (cc=131 and ll>=155 and ll<167)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="0111")) then
	if ((cc=69 and ll=137) or (cc=70 and ll=137) or (cc=71 and ll>=137 and ll<139) or (cc=72 and ll=138) or (cc=73 and ll=138) or (cc=74 and ll=139) or (cc=75 and ll=139) or (cc=76 and ll>=139 and ll<141) or (cc=77 and ll=140) or (cc=78 and ll>=140 and ll<142) or (cc=79 and ll=141) or (cc=80 and ll>=141 and ll<143) or (cc=81 and ll>=142 and ll<144) or (cc=82 and ll>=142 and ll<144) or (cc=83 and ll>=142 and ll<145) or (cc=84 and ll>=143 and ll<145) or (cc=85 and ll>=143 and ll<145) or (cc=86 and ll>=142 and ll<146) or (cc=87 and ll>=142 and ll<146) or (cc=88 and ll>=142 and ll<147) or (cc=89 and ll>=143 and ll<147) or (cc=90 and ll>=143 and ll<148) or (cc=91 and ll>=144 and ll<149) or (cc=92 and ll>=144 and ll<149) or (cc=93 and ll>=145 and ll<150) or (cc=94 and ll>=145 and ll<150) or (cc=95 and ll>=145 and ll<151) or (cc=96 and ll>=146 and ll<151) or (cc=97 and ll>=146 and ll<152) or (cc=98 and ll>=147 and ll<152) or (cc=99 and ll>=147 and ll<152) or (cc=100 and ll>=147 and ll<153) or (cc=101 and ll>=148 and ll<154) or (cc=102 and ll>=148 and ll<155) or (cc=103 and ll>=149 and ll<155) or (cc=104 and ll>=149 and ll<155) or (cc=105 and ll>=149 and ll<156) or (cc=106 and ll>=150 and ll<156) or (cc=107 and ll>=149 and ll<157) or (cc=108 and ll>=149 and ll<157) or (cc=109 and ll>=149 and ll<157) or (cc=110 and ll>=150 and ll<158) or (cc=111 and ll>=150 and ll<158) or (cc=112 and ll>=150 and ll<160) or (cc=113 and ll>=151 and ll<160) or (cc=114 and ll>=151 and ll<161) or (cc=115 and ll>=152 and ll<161) or (cc=116 and ll>=152 and ll<161) or (cc=117 and ll>=152 and ll<162) or (cc=118 and ll>=153 and ll<162) or (cc=119 and ll>=153 and ll<163) or (cc=120 and ll>=154 and ll<163) or (cc=121 and ll>=154 and ll<163) or (cc=122 and ll>=155 and ll<164) or (cc=123 and ll>=155 and ll<165) or (cc=124 and ll>=155 and ll<166) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=156 and ll<167) or (cc=127 and ll>=157 and ll<167) or (cc=128 and ll>=157 and ll<168) or (cc=129 and ll>=156 and ll<168) or (cc=130 and ll>=156 and ll<168) or (cc=131 and ll>=156 and ll<166)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="1000")) then
	if ((cc=71 and ll>=125 and ll<127) or (cc=72 and ll=126) or (cc=73 and ll>=126 and ll<128) or (cc=74 and ll=127) or (cc=75 and ll=128) or (cc=76 and ll=129) or (cc=77 and ll=129) or (cc=78 and ll=130) or (cc=79 and ll>=130 and ll<132) or (cc=80 and ll=131) or (cc=81 and ll>=132 and ll<134) or (cc=82 and ll>=132 and ll<135) or (cc=83 and ll>=133 and ll<135) or (cc=84 and ll>=133 and ll<136) or (cc=85 and ll>=134 and ll<137) or (cc=86 and ll>=135 and ll<137) or (cc=87 and ll>=133 and ll<138) or (cc=88 and ll>=134 and ll<138) or (cc=89 and ll>=135 and ll<139) or (cc=90 and ll>=135 and ll<140) or (cc=91 and ll>=136 and ll<142) or (cc=92 and ll>=137 and ll<142) or (cc=93 and ll>=137 and ll<143) or (cc=94 and ll>=138 and ll<143) or (cc=95 and ll>=139 and ll<144) or (cc=96 and ll>=139 and ll<145) or (cc=97 and ll>=140 and ll<145) or (cc=98 and ll>=140 and ll<146) or (cc=99 and ll>=141 and ll<147) or (cc=100 and ll>=142 and ll<147) or (cc=101 and ll>=142 and ll<148) or (cc=102 and ll>=143 and ll<150) or (cc=103 and ll>=144 and ll<150) or (cc=104 and ll>=144 and ll<151) or (cc=105 and ll>=145 and ll<152) or (cc=106 and ll>=146 and ll<152) or (cc=107 and ll>=146 and ll<153) or (cc=108 and ll>=145 and ll<153) or (cc=109 and ll>=146 and ll<154) or (cc=110 and ll>=146 and ll<155) or (cc=111 and ll>=147 and ll<155) or (cc=112 and ll>=147 and ll<157) or (cc=113 and ll>=148 and ll<158) or (cc=114 and ll>=149 and ll<158) or (cc=115 and ll>=149 and ll<159) or (cc=116 and ll>=150 and ll<160) or (cc=117 and ll>=150 and ll<160) or (cc=118 and ll>=151 and ll<161) or (cc=119 and ll>=152 and ll<161) or (cc=120 and ll>=153 and ll<162) or (cc=121 and ll>=153 and ll<163) or (cc=122 and ll>=154 and ll<165) or (cc=123 and ll>=154 and ll<165) or (cc=124 and ll>=155 and ll<166) or (cc=125 and ll>=156 and ll<166) or (cc=126 and ll>=156 and ll<167) or (cc=127 and ll>=157 and ll<168) or (cc=128 and ll>=157 and ll<168) or (cc=129 and ll>=156 and ll<169) or (cc=130 and ll>=157 and ll<169) or (cc=131 and ll>=157 and ll<166) or (cc=132 and ll=158)) then grbp<="101";
	end if;

elsif ((PT4 ="0100" and PT5 ="1001")) then
	if ((cc=73 and ll=114) or (cc=74 and ll=115) or (cc=75 and ll=116) or (cc=76 and ll>=116 and ll<118) or (cc=77 and ll=118) or (cc=78 and ll=119) or (cc=79 and ll>=119 and ll<121) or (cc=80 and ll>=120 and ll<122) or (cc=81 and ll=121) or (cc=82 and ll>=122 and ll<124) or (cc=83 and ll>=123 and ll<125) or (cc=84 and ll>=124 and ll<126) or (cc=85 and ll>=125 and ll<127) or (cc=86 and ll>=125 and ll<128) or (cc=87 and ll>=126 and ll<129) or (cc=88 and ll>=126 and ll<130) or (cc=89 and ll>=126 and ll<130) or (cc=90 and ll>=127 and ll<132) or (cc=91 and ll>=128 and ll<133) or (cc=92 and ll>=128 and ll<133) or (cc=93 and ll>=130 and ll<135) or (cc=94 and ll>=130 and ll<136) or (cc=95 and ll>=131 and ll<137) or (cc=96 and ll>=132 and ll<138) or (cc=97 and ll>=133 and ll<139) or (cc=98 and ll>=134 and ll<139) or (cc=99 and ll>=135 and ll<141) or (cc=100 and ll>=136 and ll<141) or (cc=101 and ll>=136 and ll<142) or (cc=102 and ll>=137 and ll<144) or (cc=103 and ll>=138 and ll<145) or (cc=104 and ll>=139 and ll<146) or (cc=105 and ll>=140 and ll<147) or (cc=106 and ll>=141 and ll<148) or (cc=107 and ll>=142 and ll<149) or (cc=108 and ll>=142 and ll<150) or (cc=109 and ll>=141 and ll<150) or (cc=110 and ll>=142 and ll<151) or (cc=111 and ll>=143 and ll<152) or (cc=112 and ll>=144 and ll<154) or (cc=113 and ll>=145 and ll<155) or (cc=114 and ll>=146 and ll<156) or (cc=115 and ll>=147 and ll<157) or (cc=116 and ll>=147 and ll<158) or (cc=117 and ll>=148 and ll<159) or (cc=118 and ll>=149 and ll<159) or (cc=119 and ll>=150 and ll<160) or (cc=120 and ll>=151 and ll<161) or (cc=121 and ll>=152 and ll<162) or (cc=122 and ll>=153 and ll<164) or (cc=123 and ll>=154 and ll<165) or (cc=124 and ll>=154 and ll<166) or (cc=125 and ll>=156 and ll<167) or (cc=126 and ll>=156 and ll<168) or (cc=127 and ll>=157 and ll<168) or (cc=128 and ll>=158 and ll<169) or (cc=129 and ll>=157 and ll<170) or (cc=130 and ll>=158 and ll<169) or (cc=131 and ll>=159 and ll<164) or (cc=132 and ll=159)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0000")) then
	if ((cc=76 and ll>=103 and ll<105) or (cc=77 and ll=105) or (cc=78 and ll=106) or (cc=79 and ll>=107 and ll<109) or (cc=80 and ll>=108 and ll<110) or (cc=81 and ll>=109 and ll<111) or (cc=82 and ll>=110 and ll<112) or (cc=83 and ll=112) or (cc=84 and ll=113) or (cc=85 and ll>=114 and ll<117) or (cc=86 and ll>=115 and ll<118) or (cc=87 and ll>=116 and ll<119) or (cc=88 and ll>=117 and ll<120) or (cc=89 and ll>=118 and ll<121) or (cc=90 and ll>=118 and ll<123) or (cc=91 and ll>=119 and ll<124) or (cc=92 and ll>=120 and ll<125) or (cc=93 and ll>=121 and ll<126) or (cc=94 and ll>=122 and ll<128) or (cc=95 and ll>=123 and ll<129) or (cc=96 and ll>=124 and ll<130) or (cc=97 and ll>=126 and ll<131) or (cc=98 and ll>=126 and ll<133) or (cc=99 and ll>=127 and ll<134) or (cc=100 and ll>=129 and ll<135) or (cc=101 and ll>=130 and ll<136) or (cc=102 and ll>=131 and ll<137) or (cc=103 and ll>=132 and ll<140) or (cc=104 and ll>=133 and ll<141) or (cc=105 and ll>=134 and ll<142) or (cc=106 and ll>=135 and ll<143) or (cc=107 and ll>=137 and ll<144) or (cc=108 and ll>=138 and ll<145) or (cc=109 and ll>=139 and ll<147) or (cc=110 and ll>=138 and ll<148) or (cc=111 and ll>=139 and ll<149) or (cc=112 and ll>=140 and ll<150) or (cc=113 and ll>=141 and ll<152) or (cc=114 and ll>=143 and ll<154) or (cc=115 and ll>=144 and ll<155) or (cc=116 and ll>=145 and ll<156) or (cc=117 and ll>=146 and ll<157) or (cc=118 and ll>=147 and ll<158) or (cc=119 and ll>=148 and ll<159) or (cc=120 and ll>=150 and ll<160) or (cc=121 and ll>=151 and ll<161) or (cc=122 and ll>=152 and ll<164) or (cc=123 and ll>=153 and ll<165) or (cc=124 and ll>=154 and ll<166) or (cc=125 and ll>=155 and ll<167) or (cc=126 and ll>=156 and ll<168) or (cc=127 and ll>=158 and ll<169) or (cc=128 and ll>=159 and ll<170) or (cc=129 and ll>=160 and ll<171) or (cc=130 and ll>=158 and ll<169) or (cc=131 and ll>=160 and ll<165) or (cc=132 and ll=161)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0001")) then
	if ((cc=79 and ll>=93 and ll<95) or (cc=80 and ll>=95 and ll<97) or (cc=81 and ll>=96 and ll<98) or (cc=82 and ll>=97 and ll<100) or (cc=83 and ll>=99 and ll<101) or (cc=84 and ll>=100 and ll<103) or (cc=85 and ll>=102 and ll<104) or (cc=86 and ll>=103 and ll<105) or (cc=87 and ll>=105 and ll<108) or (cc=88 and ll>=106 and ll<109) or (cc=89 and ll>=108 and ll<111) or (cc=90 and ll>=109 and ll<112) or (cc=91 and ll>=110 and ll<114) or (cc=92 and ll>=112 and ll<115) or (cc=93 and ll>=111 and ll<117) or (cc=94 and ll>=112 and ll<118) or (cc=95 and ll>=114 and ll<120) or (cc=96 and ll>=115 and ll<122) or (cc=97 and ll>=117 and ll<123) or (cc=98 and ll>=118 and ll<125) or (cc=99 and ll>=120 and ll<126) or (cc=100 and ll>=121 and ll<128) or (cc=101 and ll>=123 and ll<129) or (cc=102 and ll>=124 and ll<130) or (cc=103 and ll>=126 and ll<132) or (cc=104 and ll>=127 and ll<133) or (cc=105 and ll>=129 and ll<137) or (cc=106 and ll>=130 and ll<138) or (cc=107 and ll>=131 and ll<139) or (cc=108 and ll>=133 and ll<141) or (cc=109 and ll>=134 and ll<142) or (cc=110 and ll>=136 and ll<144) or (cc=111 and ll>=135 and ll<145) or (cc=112 and ll>=136 and ll<146) or (cc=113 and ll>=137 and ll<149) or (cc=114 and ll>=139 and ll<151) or (cc=115 and ll>=140 and ll<152) or (cc=116 and ll>=142 and ll<153) or (cc=117 and ll>=143 and ll<155) or (cc=118 and ll>=144 and ll<156) or (cc=119 and ll>=146 and ll<158) or (cc=120 and ll>=147 and ll<159) or (cc=121 and ll>=149 and ll<161) or (cc=122 and ll>=150 and ll<163) or (cc=123 and ll>=151 and ll<164) or (cc=124 and ll>=153 and ll<166) or (cc=125 and ll>=154 and ll<167) or (cc=126 and ll>=156 and ll<169) or (cc=127 and ll>=157 and ll<170) or (cc=128 and ll>=159 and ll<172) or (cc=129 and ll>=160 and ll<171) or (cc=130 and ll>=159 and ll<169) or (cc=131 and ll>=161 and ll<165) or (cc=132 and ll=162)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0010")) then
	if ((cc=82 and ll=84) or (cc=83 and ll=85) or (cc=84 and ll>=86 and ll<88) or (cc=85 and ll>=88 and ll<90) or (cc=86 and ll>=90 and ll<92) or (cc=87 and ll>=91 and ll<94) or (cc=88 and ll>=93 and ll<96) or (cc=89 and ll>=95 and ll<97) or (cc=90 and ll>=97 and ll<100) or (cc=91 and ll>=99 and ll<102) or (cc=92 and ll>=101 and ll<104) or (cc=93 and ll>=102 and ll<106) or (cc=94 and ll>=104 and ll<108) or (cc=95 and ll>=105 and ll<109) or (cc=96 and ll>=105 and ll<111) or (cc=97 and ll>=107 and ll<113) or (cc=98 and ll>=109 and ll<116) or (cc=99 and ll>=111 and ll<118) or (cc=100 and ll>=112 and ll<120) or (cc=101 and ll>=114 and ll<121) or (cc=102 and ll>=116 and ll<123) or (cc=103 and ll>=117 and ll<125) or (cc=104 and ll>=119 and ll<127) or (cc=105 and ll>=121 and ll<129) or (cc=106 and ll>=123 and ll<132) or (cc=107 and ll>=125 and ll<133) or (cc=108 and ll>=127 and ll<135) or (cc=109 and ll>=128 and ll<137) or (cc=110 and ll>=130 and ll<139) or (cc=111 and ll>=132 and ll<141) or (cc=112 and ll>=134 and ll<143) or (cc=113 and ll>=132 and ll<144) or (cc=114 and ll>=134 and ll<147) or (cc=115 and ll>=136 and ll<149) or (cc=116 and ll>=138 and ll<151) or (cc=117 and ll>=140 and ll<153) or (cc=118 and ll>=142 and ll<155) or (cc=119 and ll>=144 and ll<156) or (cc=120 and ll>=145 and ll<158) or (cc=121 and ll>=147 and ll<160) or (cc=122 and ll>=149 and ll<163) or (cc=123 and ll>=150 and ll<165) or (cc=124 and ll>=152 and ll<167) or (cc=125 and ll>=154 and ll<168) or (cc=126 and ll>=156 and ll<170) or (cc=127 and ll>=158 and ll<172) or (cc=128 and ll>=160 and ll<173) or (cc=129 and ll>=161 and ll<170) or (cc=130 and ll>=160 and ll<167) or (cc=131 and ll>=162 and ll<166)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0011")) then
	if ((cc=87 and ll>=76 and ll<78) or (cc=88 and ll>=78 and ll<80) or (cc=89 and ll>=80 and ll<83) or (cc=90 and ll>=82 and ll<85) or (cc=91 and ll>=85 and ll<87) or (cc=92 and ll>=87 and ll<89) or (cc=93 and ll>=89 and ll<91) or (cc=94 and ll>=91 and ll<95) or (cc=95 and ll>=93 and ll<97) or (cc=96 and ll>=96 and ll<99) or (cc=97 and ll>=98 and ll<102) or (cc=98 and ll>=100 and ll<104) or (cc=99 and ll>=99 and ll<106) or (cc=100 and ll>=101 and ll<108) or (cc=101 and ll>=103 and ll<112) or (cc=102 and ll>=105 and ll<114) or (cc=103 and ll>=108 and ll<116) or (cc=104 and ll>=110 and ll<119) or (cc=105 and ll>=112 and ll<121) or (cc=106 and ll>=114 and ll<123) or (cc=107 and ll>=116 and ll<125) or (cc=108 and ll>=119 and ll<129) or (cc=109 and ll>=121 and ll<131) or (cc=110 and ll>=123 and ll<133) or (cc=111 and ll>=125 and ll<136) or (cc=112 and ll>=128 and ll<138) or (cc=113 and ll>=130 and ll<140) or (cc=114 and ll>=130 and ll<142) or (cc=115 and ll>=131 and ll<146) or (cc=116 and ll>=134 and ll<148) or (cc=117 and ll>=136 and ll<150) or (cc=118 and ll>=138 and ll<153) or (cc=119 and ll>=140 and ll<155) or (cc=120 and ll>=143 and ll<157) or (cc=121 and ll>=145 and ll<159) or (cc=122 and ll>=147 and ll<163) or (cc=123 and ll>=149 and ll<165) or (cc=124 and ll>=151 and ll<167) or (cc=125 and ll>=154 and ll<169) or (cc=126 and ll>=156 and ll<171) or (cc=127 and ll>=158 and ll<173) or (cc=128 and ll>=160 and ll<173) or (cc=129 and ll>=162 and ll<171) or (cc=130 and ll>=161 and ll<169) or (cc=131 and ll>=163 and ll<167)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0100")) then
	if ((cc=91 and ll=68) or (cc=92 and ll>=69 and ll<72) or (cc=93 and ll>=72 and ll<75) or (cc=94 and ll>=75 and ll<77) or (cc=95 and ll>=77 and ll<80) or (cc=96 and ll>=80 and ll<83) or (cc=97 and ll>=83 and ll<87) or (cc=98 and ll>=85 and ll<90) or (cc=99 and ll>=88 and ll<93) or (cc=100 and ll>=91 and ll<95) or (cc=101 and ll>=94 and ll<98) or (cc=102 and ll>=93 and ll<101) or (cc=103 and ll>=96 and ll<106) or (cc=104 and ll>=98 and ll<108) or (cc=105 and ll>=101 and ll<111) or (cc=106 and ll>=104 and ll<114) or (cc=107 and ll>=106 and ll<116) or (cc=108 and ll>=110 and ll<119) or (cc=109 and ll>=112 and ll<122) or (cc=110 and ll>=114 and ll<126) or (cc=111 and ll>=118 and ll<129) or (cc=112 and ll>=120 and ll<131) or (cc=113 and ll>=123 and ll<135) or (cc=114 and ll>=126 and ll<137) or (cc=115 and ll>=128 and ll<139) or (cc=116 and ll>=128 and ll<144) or (cc=117 and ll>=130 and ll<147) or (cc=118 and ll>=133 and ll<150) or (cc=119 and ll>=136 and ll<152) or (cc=120 and ll>=138 and ll<155) or (cc=121 and ll>=142 and ll<158) or (cc=122 and ll>=144 and ll<162) or (cc=123 and ll>=147 and ll<165) or (cc=124 and ll>=150 and ll<168) or (cc=125 and ll>=152 and ll<170) or (cc=126 and ll>=155 and ll<173) or (cc=127 and ll>=158 and ll<174) or (cc=128 and ll>=161 and ll<172) or (cc=129 and ll>=162 and ll<171) or (cc=130 and ll>=163 and ll<168) or (cc=131 and ll>=165 and ll<167)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0101")) then
	if ((cc=96 and ll=62) or (cc=97 and ll>=62 and ll<66) or (cc=98 and ll>=66 and ll<69) or (cc=99 and ll>=69 and ll<73) or (cc=100 and ll>=73 and ll<76) or (cc=101 and ll>=76 and ll<82) or (cc=102 and ll>=80 and ll<85) or (cc=103 and ll>=83 and ll<89) or (cc=104 and ll>=87 and ll<92) or (cc=105 and ll>=89 and ll<96) or (cc=106 and ll>=90 and ll<102) or (cc=107 and ll>=93 and ll<104) or (cc=108 and ll>=97 and ll<108) or (cc=109 and ll>=100 and ll<111) or (cc=110 and ll>=104 and ll<115) or (cc=111 and ll>=107 and ll<118) or (cc=112 and ll>=110 and ll<124) or (cc=113 and ll>=113 and ll<127) or (cc=114 and ll>=117 and ll<131) or (cc=115 and ll>=120 and ll<134) or (cc=116 and ll>=124 and ll<137) or (cc=117 and ll>=126 and ll<143) or (cc=118 and ll>=127 and ll<147) or (cc=119 and ll>=130 and ll<150) or (cc=120 and ll>=134 and ll<153) or (cc=121 and ll>=137 and ll<156) or (cc=122 and ll>=141 and ll<162) or (cc=123 and ll>=144 and ll<165) or (cc=124 and ll>=148 and ll<169) or (cc=125 and ll>=151 and ll<172) or (cc=126 and ll>=155 and ll<174) or (cc=127 and ll>=158 and ll<173) or (cc=128 and ll>=161 and ll<172) or (cc=129 and ll>=163 and ll<170) or (cc=130 and ll>=164 and ll<169) or (cc=131 and ll=167)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0110")) then
	if ((cc=102 and ll>=56 and ll<61) or (cc=103 and ll>=61 and ll<65) or (cc=104 and ll>=65 and ll<70) or (cc=105 and ll>=70 and ll<74) or (cc=106 and ll>=74 and ll<81) or (cc=107 and ll>=78 and ll<86) or (cc=108 and ll>=83 and ll<89) or (cc=109 and ll>=85 and ll<94) or (cc=110 and ll>=87 and ll<101) or (cc=111 and ll>=91 and ll<105) or (cc=112 and ll>=95 and ll<110) or (cc=113 and ll>=100 and ll<114) or (cc=114 and ll>=104 and ll<121) or (cc=115 and ll>=109 and ll<126) or (cc=116 and ll>=114 and ll<130) or (cc=117 and ll>=118 and ll<135) or (cc=118 and ll>=123 and ll<142) or (cc=119 and ll>=125 and ll<146) or (cc=120 and ll>=126 and ll<150) or (cc=121 and ll>=131 and ll<154) or (cc=122 and ll>=136 and ll<161) or (cc=123 and ll>=139 and ll<166) or (cc=124 and ll>=144 and ll<170) or (cc=125 and ll>=148 and ll<174) or (cc=126 and ll>=153 and ll<174) or (cc=127 and ll>=157 and ll<173) or (cc=128 and ll>=162 and ll<171) or (cc=129 and ll>=164 and ll<170) or (cc=130 and ll>=166 and ll<169)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="0111")) then
	if ((cc=107 and ll>=52 and ll<55) or (cc=108 and ll>=55 and ll<60) or (cc=109 and ll>=60 and ll<67) or (cc=110 and ll>=67 and ll<76) or (cc=111 and ll>=73 and ll<82) or (cc=112 and ll>=78 and ll<88) or (cc=113 and ll>=82 and ll<97) or (cc=114 and ll>=84 and ll<104) or (cc=115 and ll>=90 and ll<109) or (cc=116 and ll>=97 and ll<118) or (cc=117 and ll>=102 and ll<125) or (cc=118 and ll>=109 and ll<131) or (cc=119 and ll>=115 and ll<140) or (cc=120 and ll>=120 and ll<146) or (cc=121 and ll>=124 and ll<152) or (cc=122 and ll>=126 and ll<162) or (cc=123 and ll>=132 and ll<167) or (cc=124 and ll>=139 and ll<173) or (cc=125 and ll>=145 and ll<174) or (cc=126 and ll>=151 and ll<173) or (cc=127 and ll>=157 and ll<172) or (cc=128 and ll>=163 and ll<172) or (cc=129 and ll>=165 and ll<171) or (cc=130 and ll>=169 and ll<171)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="1000")) then
	if ((cc=113 and ll>=49 and ll<54) or (cc=114 and ll>=54 and ll<64) or (cc=115 and ll>=64 and ll<78) or (cc=116 and ll>=73 and ll<87) or (cc=117 and ll>=80 and ll<101) or (cc=118 and ll>=82 and ll<115) or (cc=119 and ll>=91 and ll<125) or (cc=120 and ll>=101 and ll<138) or (cc=121 and ll>=110 and ll<147) or (cc=122 and ll>=119 and ll<161) or (cc=123 and ll>=123 and ll<170) or (cc=124 and ll>=128 and ll<174) or (cc=125 and ll>=137 and ll<173) or (cc=126 and ll>=146 and ll<173) or (cc=127 and ll>=155 and ll<172) or (cc=128 and ll>=165 and ll<172) or (cc=129 and ll>=166 and ll<171)) then grbp<="101";
	end if;

elsif ((PT4 ="0101" and PT5 ="1001")) then
	if ((cc=119 and ll>=47 and ll<70) or (cc=120 and ll>=61 and ll<97) or (cc=121 and ll>=78 and ll<125) or (cc=122 and ll>=79 and ll<161) or (cc=123 and ll>=97 and ll<173) or (cc=124 and ll>=115 and ll<173) or (cc=125 and ll>=123 and ll<173) or (cc=126 and ll>=133 and ll<173) or (cc=127 and ll>=152 and ll<173) or (cc=128 and ll>=166 and ll<172) or (cc=129 and ll>=169 and ll<172)) then grbp<="101";
	end if;


end if;

	IF CC >85 and cc<90 AND ((LL <330 AND LL > 320) or (ll<380 and ll>370)) THEN GRBP <= "111";
	END IF;

	IF CC >160 and cc<165 AND ((LL <330 AND LL > 320) or (ll<380 and ll>370)) THEN GRBP <= "111";
	END IF;

if PT0="0000" then
	if (cc>30 and cc<46 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>30 and cc<36 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>40 and cc<46 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>30 and cc<46 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT0="0001" then
	if (cc>35 and cc<41 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT0="0010" then
	if (cc>30 and cc<46 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>40 and cc<46 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>30 and cc<46 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>30 and cc<36 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>30 and cc<46 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

if PT1="0000" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>55 and cc<60 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>66 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0001" then
	if (cc>60 and cc<66 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0010" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<61 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0011" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0100" then
	if (cc>55 and cc<61 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0101" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>55 and cc<61 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0110" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>55 and cc<61 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="0111" then
	if (cc>55 and cc<61 and ll>310 and ll<319) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="1000" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>55 and cc<61 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT1="1001" then
	if (cc>55 and cc<71 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>55 and cc<61 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>65 and cc<71 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>55 and cc<71 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

if PT2="0000" then
	if (cc>105 and cc<121 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>105 and cc<110 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>116 and cc<121 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT2="0001" then
	if (cc>110 and cc<116 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT2="0010" then
	if (cc>105 and cc<121 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>115 and cc<121 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>105 and cc<111 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT2="0011" then
	if (cc>105 and cc<121 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>115 and cc<121 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT2="0100" then
	if (cc>105 and cc<111 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>115 and cc<121 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT2="0101" then
	if (cc>105 and cc<121 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>105 and cc<111 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>115 and cc<121 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>105 and cc<121 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

if PT3="0000" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0001" then
	if (cc>135 and cc<141 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0010" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0011" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0100" then
	if (cc>130 and cc<136 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0101" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0110" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="0111" then
	if (cc>130 and cc<136 and ll>310 and ll<319) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="1000" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT3="1001" then
	if (cc>130 and cc<146 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>130 and cc<136 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>140 and cc<146 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>130 and cc<146 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

if PT4="0000" then
	if (cc>180 and cc<196 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>180 and cc<186 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>190 and cc<196 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT4="0001" then
	if (cc>185 and cc<191 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT4="0010" then
	if (cc>180 and cc<196 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>190 and cc<196 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>180 and cc<186 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT4="0011" then
	if (cc>180 and cc<196 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>190 and cc<196 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT4="0100" then
	if (cc>180 and cc<186 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>190 and cc<196 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT4="0101" then
	if (cc>180 and cc<196 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>180 and cc<186 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>190 and cc<196 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>180 and cc<196 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

if PT5="0000" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>205 and cc<210 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>216 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0001" then
	if (cc>210 and cc<216 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0010" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<211 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0011" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0100" then
	if (cc>205 and cc<211 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0101" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>205 and cc<211 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0110" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>205 and cc<211 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>342 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="0111" then
	if (cc>205 and cc<211 and ll>310 and ll<319) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="1000" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>205 and cc<211 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;
if PT5="1001" then
	if (cc>205 and cc<221 and ll>310 and ll<327) then grbp<="010";
	end if;
	if (cc>205 and cc<211 and ll>310 and ll<359) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>342 and ll<359) then grbp<="010";
	end if;
	if (cc>215 and cc<221 and ll>310 and ll<391) then grbp<="010";
	end if;
	if (cc>205 and cc<221 and ll>374 and ll<391) then grbp<="010";
	end if;
end if;

end if;
-------------------------------mode="101"--------------------wave--------------------
if mode="101" then
cci<=to_integer(unsigned(cc));

if (cci>26 and cci<226) then
	if (tri='1' and ll=tri_ind(cci-25)+90) then grbp<="100";
	end if;
	if (squ='1' and ll=squ_ind(cci-25)+90) then grbp<="010";
    end if;
	if (sin='1' and  ll=sin_id(cci-25)+90) then grbp<="011";
    end if;
end if;	

if cc>26 and cc<226 and ll>89 and ll<291 then
if cc=rrll+26 then
    grbp<="101";
end if;

if ll=190 then
    grbp<="101";
end if;
end if;

if cc=26 and ll>89 and ll<291 then
    grbp<="111";
end if;

--------------------------xscal--------begin----40-55-56-71--295-335----------

	if (cc=41 and ll=297) then grbp<="010";
	end if;
	if (ll=297 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=297 and cc>=50 and cc<54) then grbp<="010";
	end if;
	if (cc=41 and ll=298) then grbp<="010";
	end if;
	if (ll=298 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=298 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=299 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=299 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=300 and cc>=42 and cc<45) then grbp<="010";
	end if;
	if (ll=300 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=301 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=301 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=302 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=302 and cc>=49 and cc<52) then grbp<="010";
	end if;
	if (ll=303 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=303 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=304 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=304 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=305 and cc>=43 and cc<47) then grbp<="010";
	end if;
	if (ll=305 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=306 and cc>=43 and cc<47) then grbp<="010";
	end if;
	if (ll=306 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=307 and cc>=43 and cc<51) then grbp<="010";
	end if;
	if (ll=308 and cc>=44 and cc<51) then grbp<="010";
	end if;
	if (ll=309 and cc>=44 and cc<51) then grbp<="010";
	end if;
	if (ll=310 and cc>=44 and cc<51) then grbp<="010";
	end if;
	if (ll=311 and cc>=44 and cc<50) then grbp<="010";
	end if;
	if (ll=312 and cc>=45 and cc<50) then grbp<="010";
	end if;
	if (ll=313 and cc>=45 and cc<50) then grbp<="010";
	end if;
	if (ll=314 and cc>=45 and cc<50) then grbp<="010";
	end if;
	if (ll=315 and cc>=45 and cc<50) then grbp<="010";
	end if;
	if (ll=316 and cc>=44 and cc<50) then grbp<="010";
	end if;
	if (ll=317 and cc>=44 and cc<50) then grbp<="010";
	end if;
	if (ll=318 and cc>=44 and cc<50) then grbp<="010";
	end if;
	if (ll=319 and cc>=44 and cc<51) then grbp<="010";
	end if;
	if (ll=320 and cc>=43 and cc<51) then grbp<="010";
	end if;
	if (ll=321 and cc>=43 and cc<51) then grbp<="010";
	end if;
	if (ll=322 and cc>=43 and cc<47) then grbp<="010";
	end if;
	if (ll=322 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=323 and cc>=43 and cc<47) then grbp<="010";
	end if;
	if (ll=323 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=324 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=324 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=325 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=325 and cc>=48 and cc<52) then grbp<="010";
	end if;
	if (ll=326 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=326 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=327 and cc>=42 and cc<46) then grbp<="010";
	end if;
	if (ll=327 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=328 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=328 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=329 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=329 and cc>=49 and cc<53) then grbp<="010";
	end if;
	if (ll=330 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=330 and cc>=50 and cc<54) then grbp<="010";
	end if;
	if (cc=41 and ll=331) then grbp<="010";
	end if;
	if (ll=331 and cc>=41 and cc<45) then grbp<="010";
	end if;
	if (ll=331 and cc>=50 and cc<54) then grbp<="010";
	end if;



if sc=1 then
	if (cc>61 and cc<67 and ll>295 and ll<336) then grbp<="010";
	end if;
end if;
if sc=2 then
	if (cc>56 and cc<72 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>66 and cc<72 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>56 and cc<72 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>56 and cc<62 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>56 and cc<72 and ll>327 and ll<336) then grbp<="010";
	end if;
end if;
if sc=4 then
	if (cc>56 and cc<62 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>56 and cc<72 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>66 and cc<72 and ll>295 and ll<336) then grbp<="010";
	end if;
end if;
if sc=8 then
	if (cc>56 and cc<72 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>56 and cc<62 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>56 and cc<72 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>66 and cc<72 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>56 and cc<72 and ll>327 and ll<336) then grbp<="010";
	end if;
end if;

---------------------------xscal-------end-----------------

---------------------------T-----begin----225-190----------

if sc=1 then

	if (cc>219 and cc<222 and ll>191 and ll<200) then grbp<="011";
	end if;
	if (cc>219 and cc<225 and ll>197 and ll<200) then grbp<="011";
	end if;
	if (cc>222 and cc<225 and ll>191 and ll<206) then grbp<="011";
	end if;
	
end if;

if sc=2 then
    
	if (cc>219 and cc<225 and ll>191 and ll<195) then grbp<="011";
	end if;
	if (cc>222 and cc<225 and ll>191 and ll<200) then grbp<="011";
	end if;
	if (cc>219 and cc<225 and ll>197 and ll<200) then grbp<="011";
	end if;
	if (cc>219 and cc<222 and ll>197 and ll<206) then grbp<="011";
	end if;
	if (cc>219 and cc<225 and ll>202 and ll<206) then grbp<="011";
	end if;

end if;

if sc=4 then

	if (cc=222 and ll>191 and ll<206) then grbp<="011";
	end if;
	
end if;

if sc=1 or sc=2 or sc=4 then

    if (cc=228 and ll=195) then grbp<="011";
	end if;
	if (cc=225 and ll=196) then grbp<="011";
	end if;
	if (cc=228 and ll=196) then grbp<="011";
	end if;
	if (cc=225 and ll=197) then grbp<="011";
	end if;
	if (cc=228 and ll=197) then grbp<="011";
	end if;
	if (cc=225 and ll=198) then grbp<="011";
	end if;
	if (cc=228 and ll=198) then grbp<="011";
	end if;
	if (cc=225 and ll=199) then grbp<="011";
	end if;
	if (cc=228 and ll=199) then grbp<="011";
	end if;
	if (cc=225 and ll=200) then grbp<="011";
	end if;
	if (cc=228 and ll=200) then grbp<="011";
	end if;
	if (cc=225 and ll=201) then grbp<="011";
	end if;
	if (cc=228 and ll=201) then grbp<="011";
	end if;
	if (cc=225 and ll=202) then grbp<="011";
	end if;
	if (ll=202 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (cc=225 and ll=203) then grbp<="011";
	end if;
	if (ll=203 and cc>=225 and cc<230) then grbp<="011";
	end if;
	if (ll=204 and cc>=225 and cc<228) then grbp<="011";
	end if;
	if (cc=225 and ll=205) then grbp<="011";
	end if;
	if (cc=225 and ll=206) then grbp<="011";
	end if;

end if;

if sc=8 then

	if (cc>207 and cc<213 and ll>191 and ll<195) then grbp<="011";
	end if;
	if (cc>207 and cc<210 and ll>191 and ll<200) then grbp<="011";
	end if;
	if (cc>207 and cc<213 and ll>197 and ll<200) then grbp<="011";
	end if;
	if (cc>210 and cc<213 and ll>197 and ll<206) then grbp<="011";
	end if;
	if (cc>207 and cc<213 and ll>202 and ll<206) then grbp<="011";
	end if;

	if (cc>213 and cc<219 and ll>191 and ll<195) then grbp<="011";
	end if;
	if (cc>213 and cc<216 and ll>191 and ll<206) then grbp<="011";
	end if;
	if (cc>216 and cc<219 and ll>191 and ll<206) then grbp<="011";
	end if;
	if (cc>213 and cc<219 and ll>202 and ll<206) then grbp<="011";
	end if;

	if (cc>219 and cc<225 and ll>191 and ll<195) then grbp<="011";
	end if;
	if (cc>219 and cc<222 and ll>191 and ll<206) then grbp<="011";
	end if;
	if (cc>222 and cc<225 and ll>191 and ll<206) then grbp<="011";
	end if;
	if (cc>219 and cc<225 and ll>202 and ll<206) then grbp<="011";
	end if;
		
	if (cc=228 and ll=195) then grbp<="011";
	end if;
	if (cc=225 and ll=196) then grbp<="011";
	end if;
	if (cc=227 and ll=196) then grbp<="011";
	end if;
	if (ll=196 and cc>=227 and cc<229) then grbp<="011";
	end if;
	if (ll=197 and cc>=225 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=198) then grbp<="011";
	end if;
	if (ll=198 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=198 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=199) then grbp<="011";
	end if;
	if (ll=199 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=199 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=200) then grbp<="011";
	end if;
	if (ll=200 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=200 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=201) then grbp<="011";
	end if;
	if (ll=201 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=201 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=202) then grbp<="011";
	end if;
	if (ll=202 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=202 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=203) then grbp<="011";
	end if;
	if (ll=203 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=203 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=204) then grbp<="011";
	end if;
	if (ll=204 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=204 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=225 and ll=205) then grbp<="011";
	end if;
	if (ll=205 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (ll=205 and cc>=228 and cc<230) then grbp<="011";
	end if;
    
end if;

	if (cc=233 and ll=195) then grbp<="011";
	end if;
	if (cc=232 and ll=196) then grbp<="011";
	end if;
	if (ll=196 and cc>=232 and cc<235) then grbp<="011";
	end if;
	if (cc=235 and ll=196) then grbp<="011";
	end if;
	if (cc=231 and ll=197) then grbp<="011";
	end if;
	if (ll=197 and cc>=231 and cc<235) then grbp<="011";
	end if;
	if (cc=231 and ll=198) then grbp<="011";
	end if;
	if (ll=198 and cc>=231 and cc<233) then grbp<="011";
	end if;
	if (ll=199 and cc>=231 and cc<234) then grbp<="011";
	end if;
	if (ll=200 and cc>=232 and cc<235) then grbp<="011";
	end if;
	if (cc=232 and ll=201) then grbp<="011";
	end if;
	if (ll=201 and cc>=232 and cc<235) then grbp<="011";
	end if;
	if (cc=235 and ll=201) then grbp<="011";
	end if;
	if (cc=234 and ll=202) then grbp<="011";
	end if;
	if (ll=202 and cc>=234 and cc<236) then grbp<="011";
	end if;
	if (cc=234 and ll=203) then grbp<="011";
	end if;
	if (ll=203 and cc>=234 and cc<236) then grbp<="011";
	end if;
	if (ll=204 and cc>=231 and cc<235) then grbp<="011";
	end if;
	if (cc=235 and ll=204) then grbp<="011";
	end if;
	if (cc=231 and ll=205) then grbp<="011";
	end if;
	if (ll=205 and cc>=231 and cc<235) then grbp<="011";
	end if;

---------------------------T-----end------------------

-----------------------------freq-------begin----------85-100-115-130-135-150-165-180-195-210---

	if (cc>91 and cc<99 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>91 and cc<94 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>86 and cc<99 and ll>311 and ll<320) then grbp<="010";
	end if;

	if (cc>100 and cc<115 and ll>303 and ll<312) then grbp<="010";
	end if;
	if (cc>100 and cc<115 and ll>319 and ll<328) then grbp<="010";
	end if;

if f=1 then

	if (cc>120 and cc<135 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>129 and cc<135 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>120 and cc<135 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>120 and cc<126 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>120 and cc<135 and ll>327 and ll<336) then grbp<="010";
	end if;

	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>135 and cc<141 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;	
	
end if;

if f=2 then
	if (cc>120 and cc<135 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>120 and cc<126 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>120 and cc<135 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>129 and cc<135 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>120 and cc<135 and ll>327 and ll<336) then grbp<="010";
	end if;
	
	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>135 and cc<140 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>145 and cc<150 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;
    
end if;

if f=3 then
	if (cc>120 and cc<126 and ll>295 and ll<300) then grbp<="010";
	end if;
	if (cc>120 and cc<135 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>129 and cc<135 and ll>295 and ll<336) then grbp<="010";
	end if;
	
	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>135 and cc<141 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;
    
end if;


if f<4 then
    
	if (cc>150 and cc<165 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>150 and cc<155 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>160 and cc<165 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>150 and cc<165 and ll>327 and ll<336) then grbp<="010";
	end if;
		
	if (cc>165 and cc<169 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>314 and ll<316) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>315 and ll<317) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>316 and ll<318) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>317 and ll<319) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>318 and ll<320) then grbp<="010";
	end if;
	if (cc>171 and cc<174 and ll>319 and ll<321) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>320 and ll<322) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>321 and ll<323) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>322 and ll<324) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>323 and ll<325) then grbp<="010";
	end if;
	if (cc>165 and cc<169 and ll>324 and ll<326) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>325 and ll<327) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>326 and ll<328) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>327 and ll<329) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>328 and ll<330) then grbp<="010";
	end if;
	if (cc>171 and cc<174 and ll>329 and ll<331) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>330 and ll<332) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>331 and ll<333) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>332 and ll<334) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>333 and ll<335) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>334 and ll<336) then grbp<="010";
	end if;

end if;

if f>3 and f<8 then

	if (cc>120 and cc<125 and ll>295 and ll<336) then grbp<="010";
	end if;
    
end if;

if f=8 then
    
	if (cc>115 and cc<130 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>124 and cc<130 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>115 and cc<130 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>115 and cc<121 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>115 and cc<130 and ll>327 and ll<336) then grbp<="010";
	end if;
	
end if;

	if (cc>131 and cc<135 and ll>327 and ll<336) then grbp<="010";
	end if;

if f=4 or f=8 then
    
	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>135 and cc<140 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>145 and cc<150 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;
	
end if;

if f=5 then

	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>135 and cc<141 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;

end if;

if f=6 then

	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>135 and cc<141 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>327 and ll<336) then grbp<="010";
	end if;

end if;

if f=7 then
    
	if (cc>135 and cc<141 and ll>295 and ll<300) then grbp<="010";
	end if;
	if (cc>135 and cc<150 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>295 and ll<336) then grbp<="010";
	end if;
   
end if;

if f=4 or f=6 or f=8 then

	if (cc>150 and cc<165 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>150 and cc<155 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>160 and cc<165 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>150 and cc<165 and ll>327 and ll<336) then grbp<="010";
	end if;
    
end if;

if f=5 or f=7 then
   
	if (cc>150 and cc<165 and ll>295 and ll<304) then grbp<="010";
	end if;
	if (cc>150 and cc<156 and ll>295 and ll<320) then grbp<="010";
	end if;
	if (cc>150 and cc<165 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>159 and cc<165 and ll>311 and ll<336) then grbp<="010";
	end if;
	if (cc>150 and cc<165 and ll>327 and ll<336) then grbp<="010";
	end if;
	 
end if;

if f>3 then

    	if (cc>165 and cc<169 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>165 and cc<169 and ll>295 and ll<297) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>295 and ll<297) then grbp<="010";
	end if;
	if (cc>165 and cc<169 and ll>296 and ll<298) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>296 and ll<298) then grbp<="010";
	end if;
	if (cc>165 and cc<169 and ll>297 and ll<299) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>297 and ll<299) then grbp<="010";
	end if;
	if (cc>165 and cc<169 and ll>298 and ll<300) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>298 and ll<300) then grbp<="010";
	end if;
	if (cc>166 and cc<169 and ll>299 and ll<301) then grbp<="010";
	end if;
	if (cc>176 and cc<179 and ll>299 and ll<301) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>300 and ll<302) then grbp<="010";
	end if;
	if (cc>176 and cc<179 and ll>300 and ll<302) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>301 and ll<303) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>301 and ll<303) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>302 and ll<304) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>302 and ll<304) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>303 and ll<305) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>303 and ll<305) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>304 and ll<306) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>304 and ll<306) then grbp<="010";
	end if;
	if (cc>166 and cc<170 and ll>305 and ll<307) then grbp<="010";
	end if;
	if (cc>175 and cc<179 and ll>305 and ll<307) then grbp<="010";
	end if;
	if (cc>167 and cc<170 and ll>306 and ll<308) then grbp<="010";
	end if;
	if (cc>175 and cc<178 and ll>306 and ll<308) then grbp<="010";
	end if;
	if (cc>167 and cc<170 and ll>307 and ll<309) then grbp<="010";
	end if;
	if (cc>175 and cc<178 and ll>307 and ll<309) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>308 and ll<310) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>308 and ll<310) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>309 and ll<311) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>309 and ll<311) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>310 and ll<312) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>310 and ll<312) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>311 and ll<313) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>311 and ll<313) then grbp<="010";
	end if;
	if (cc>167 and cc<171 and ll>312 and ll<314) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>312 and ll<314) then grbp<="010";
	end if;
	if (cc>168 and cc<171 and ll>313 and ll<315) then grbp<="010";
	end if;
	if (cc>174 and cc<177 and ll>313 and ll<315) then grbp<="010";
	end if;
	if (cc>168 and cc<171 and ll>314 and ll<316) then grbp<="010";
	end if;
	if (cc>174 and cc<177 and ll>314 and ll<316) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>315 and ll<317) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>315 and ll<317) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>316 and ll<318) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>316 and ll<318) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>317 and ll<319) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>317 and ll<319) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>318 and ll<320) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>318 and ll<320) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>319 and ll<321) then grbp<="010";
	end if;
	if (cc>173 and cc<177 and ll>319 and ll<321) then grbp<="010";
	end if;
	if (cc>168 and cc<172 and ll>320 and ll<322) then grbp<="010";
	end if;
	if (cc>173 and cc<176 and ll>320 and ll<322) then grbp<="010";
	end if;
	if (cc>169 and cc<172 and ll>321 and ll<323) then grbp<="010";
	end if;
	if (cc>173 and cc<176 and ll>321 and ll<323) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>322 and ll<324) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>322 and ll<324) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>323 and ll<325) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>323 and ll<325) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>324 and ll<326) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>324 and ll<326) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>325 and ll<327) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>325 and ll<327) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>326 and ll<328) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>326 and ll<328) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>327 and ll<329) then grbp<="010";
	end if;
	if (cc>172 and cc<176 and ll>327 and ll<329) then grbp<="010";
	end if;
	if (cc>170 and cc<173 and ll>328 and ll<330) then grbp<="010";
	end if;
	if (cc>172 and cc<175 and ll>328 and ll<330) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>329 and ll<331) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>329 and ll<331) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>330 and ll<332) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>330 and ll<332) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>331 and ll<333) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>331 and ll<333) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>332 and ll<334) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>332 and ll<334) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>333 and ll<335) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>333 and ll<335) then grbp<="010";
	end if;
	if (cc>170 and cc<174 and ll>334 and ll<336) then grbp<="010";
	end if;
	if (cc>171 and cc<175 and ll>334 and ll<336) then grbp<="010";
	end if;
	if (cc>176 and cc<180 and ll>295 and ll<336) then grbp<="010";
	end if;

end if;


	if (cc>180 and cc<184 and ll>295 and ll<336) then grbp<="010";
	end if;
	if (cc>180 and cc<195 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>191 and cc<195 and ll>295 and ll<336) then grbp<="010";
	end if;

	if (cc>195 and cc<209 and ll>311 and ll<320) then grbp<="010";
	end if;
	if (cc>205 and cc<209 and ll>319 and ll<321) then grbp<="010";
	end if;
	if (cc>203 and cc<207 and ll>320 and ll<322) then grbp<="010";
	end if;
	if (cc>202 and cc<206 and ll>321 and ll<323) then grbp<="010";
	end if;
	if (cc>201 and cc<204 and ll>322 and ll<324) then grbp<="010";
	end if;
	if (cc>199 and cc<203 and ll>323 and ll<325) then grbp<="010";
	end if;
	if (cc>198 and cc<202 and ll>324 and ll<326) then grbp<="010";
	end if;
	if (cc>196 and cc<200 and ll>325 and ll<327) then grbp<="010";
	end if;
	if (cc>195 and cc<199 and ll>326 and ll<328) then grbp<="010";
	end if;
	if (cc>195 and cc<209 and ll>327 and ll<336) then grbp<="010";
	end if;
end if;
-------------------------------mode="110"--------------------snake---------------------

------------------------------------------mode-logo------------------------------------

if mode="000" then
    
	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=204 and ll=52) then grbp<="001";
	end if;
	if (cc=207 and ll=52) then grbp<="001";
	end if;
	if (cc=219 and ll=52) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=53) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=56 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=57 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=203 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=58 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=203 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=59 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (ll=59 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=59 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=215 and cc<219) then grbp<="001";
	end if;
	if (ll=60 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (cc=204 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (ll=61 and cc>=214 and cc<216) then grbp<="001";
	end if;
	if (cc=220 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=227 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (cc=204 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (ll=62 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=62 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=217 and ll=62) then grbp<="001";
	end if;
	if (cc=220 and ll=62) then grbp<="001";
	end if;
	if (cc=223 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (cc=205 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=63) then grbp<="001";
	end if;
	if (cc=214 and ll=63) then grbp<="001";
	end if;
	if (cc=217 and ll=63) then grbp<="001";
	end if;
	if (cc=220 and ll=63) then grbp<="001";
	end if;
	if (cc=223 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (cc=204 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=212 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=65) then grbp<="001";
	end if;
	if (cc=212 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=66) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=217 and ll=66) then grbp<="001";
	end if;
	if (cc=219 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=202 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=67 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=217 and ll=67) then grbp<="001";
	end if;
	if (cc=219 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=202 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=202 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (ll=69 and cc>=207 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=208 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=70 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=70) then grbp<="001";
	end if;
	if (cc=222 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=208 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=72 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=209 and ll=73) then grbp<="001";
	end if;
	if (cc=220 and ll=73) then grbp<="001";
	end if;
	if (cc=201 and ll=77) then grbp<="001";
	end if;
	if (ll=77 and cc>=201 and cc<229) then grbp<="001";
	end if;
	if (cc=201 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=201 and cc<229) then grbp<="001";
	end if;

	if (cc=204 and ll=51) then grbp<="011";
	end if;
	if (cc=207 and ll=51) then grbp<="011";
	end if;
	if (ll=51 and cc>=207 and cc<209) then grbp<="011";
	end if;
	if (cc=203 and ll=52) then grbp<="011";
	end if;
	if (cc=208 and ll=52) then grbp<="011";
	end if;
	if (cc=219 and ll=53) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=206 and ll=54) then grbp<="011";
	end if;
	if (cc=227 and ll=57) then grbp<="011";
	end if;
	if (cc=216 and ll=58) then grbp<="011";
	end if;
	if (cc=205 and ll=59) then grbp<="011";
	end if;
	if (cc=223 and ll=59) then grbp<="011";
	end if;
	if (cc=207 and ll=60) then grbp<="011";
	end if;
	if (cc=214 and ll=60) then grbp<="011";
	end if;
	if (cc=220 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=203 and ll=61) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=218 and ll=61) then grbp<="011";
	end if;
	if (cc=222 and ll=61) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=203 and ll=62) then grbp<="011";
	end if;
	if (cc=203 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=203 and cc<205) then grbp<="011";
	end if;
	if (cc=219 and ll=63) then grbp<="011";
	end if;
	if (cc=203 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=65) then grbp<="011";
	end if;
	if (cc=214 and ll=65) then grbp<="011";
	end if;
	if (cc=207 and ll=66) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=220 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=220 and cc<224) then grbp<="011";
	end if;
	if (ll=70 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=215 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<204) then grbp<="111";
	end if;
	if (ll=51 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=51 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=51 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=52 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=52 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=52 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=220 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=56 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=57 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=208 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=58) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=59 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=59 and cc>=224 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=224 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=61 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (cc=216 and ll=61) then grbp<="111";
	end if;
	if (cc=219 and ll=61) then grbp<="111";
	end if;
	if (cc=224 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=210 and ll=62) then grbp<="111";
	end if;
	if (cc=213 and ll=62) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (ll=62 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=62 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=62 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=221 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=63 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=64 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=65) then grbp<="111";
	end if;
	if (cc=209 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=220 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=220 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=209 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=209 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=209 and ll=70) then grbp<="111";
	end if;
	if (cc=212 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (ll=71 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=71 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=72 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<209) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (ll=73 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (cc=229 and ll=77) then grbp<="111";
	end if;
	if (cc=200 and ll=78) then grbp<="111";
	end if;
	if (cc=229 and ll=78) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="001" then
    


	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=61 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=226 and ll=52) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=229 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=204 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=223 and ll=71) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (ll=73 and cc>=223 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=65 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=226 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (cc=228 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (cc=228 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="010" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=226 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=228 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=227 and ll=65) then grbp<="011";
	end if;
	if (ll=66 and cc>=227 and cc<229) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=225 and ll=70) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="011" then
    


	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=65) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (ll=66 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=223 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=228 and ll=52) then grbp<="011";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=227 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=226 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=226 and cc<229) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=68 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=59) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=60) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=229 and ll=66) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="100" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=215 and ll=58) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=221 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (cc=213 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=61) then grbp<="001";
	end if;
	if (cc=224 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=224 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=63 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=223 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=223 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=223 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=217 and ll=52) then grbp<="011";
	end if;
	if (cc=204 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=54) then grbp<="011";
	end if;
	if (cc=225 and ll=54) then grbp<="011";
	end if;
	if (ll=54 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=205 and ll=56) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=228 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (cc=218 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=206 and ll=64) then grbp<="011";
	end if;
	if (cc=228 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=210 and ll=67) then grbp<="011";
	end if;
	if (cc=213 and ll=67) then grbp<="011";
	end if;
	if (cc=223 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=69) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=224 and ll=70) then grbp<="011";
	end if;
	if (cc=212 and ll=71) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=226 and ll=72) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=223 and ll=60) then grbp<="111";
	end if;
	if (cc=228 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (cc=226 and ll=61) then grbp<="111";
	end if;
	if (cc=229 and ll=61) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=62 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (ll=67 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=224 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=227 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=227 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;
end if;	

if mode="101" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=226 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=228 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=224 and ll=63) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=224 and ll=66) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=227 and ll=53) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=224 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=225 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=67) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=227 and ll=71) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=56 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=57 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=58 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

if mode="111" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=229 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=211 and ll=68) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=227 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=228 and ll=54) then grbp<="011";
	end if;
	if (cc=217 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=220 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=62 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=224 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=225 and ll=64) then grbp<="011";
	end if;
	if (cc=227 and ll=64) then grbp<="011";
	end if;
	if (cc=206 and ll=65) then grbp<="011";
	end if;
	if (cc=218 and ll=65) then grbp<="011";
	end if;
	if (cc=202 and ll=66) then grbp<="011";
	end if;
	if (cc=210 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=211 and ll=69) then grbp<="011";
	end if;
	if (ll=69 and cc>=211 and cc<213) then grbp<="011";
	end if;
	if (cc=222 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (cc=226 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=228 and ll=78) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=229 and ll=63) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=226 and ll=64) then grbp<="111";
	end if;
	if (cc=229 and ll=64) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=225 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=70 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;

end if;
if mode="110" then
	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (cc=217 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=205 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=227 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=210 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (cc=219 and ll=61) then grbp<="001";
	end if;
	if (cc=221 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=218 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=226 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=210 and ll=67) then grbp<="001";
	end if;
	if (cc=212 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=215 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (cc=218 and ll=70) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=71 and cc>=212 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=73) then grbp<="001";
	end if;
	if (cc=204 and ll=73) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=213 and ll=73) then grbp<="001";
	end if;
	if (cc=215 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=207 and ll=54) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=227 and ll=56) then grbp<="011";
	end if;
	if (cc=209 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=220 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=220 and cc<222) then grbp<="011";
	end if;
	if (cc=213 and ll=60) then grbp<="011";
	end if;
	if (cc=222 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=204 and ll=61) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (cc=214 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=62) then grbp<="011";
	end if;
	if (cc=218 and ll=62) then grbp<="011";
	end if;
	if (cc=221 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="011";
	end if;
	if (cc=221 and ll=63) then grbp<="011";
	end if;
	if (cc=226 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=213 and ll=65) then grbp<="011";
	end if;
	if (cc=222 and ll=65) then grbp<="011";
	end if;
	if (cc=210 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=67) then grbp<="011";
	end if;
	if (cc=224 and ll=68) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=213 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=210 and ll=71) then grbp<="011";
	end if;
	if (cc=221 and ll=71) then grbp<="011";
	end if;
	if (cc=204 and ll=72) then grbp<="011";
	end if;
	if (cc=212 and ll=72) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (cc=207 and ll=73) then grbp<="011";
	end if;
	if (cc=209 and ll=73) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;
	if (cc=218 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=223 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=51 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=54 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (cc=217 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=217 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (cc=223 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=63 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=64 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=65 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=66 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=222 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=216 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=205 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

end process;

hs<=hs1;vs<=vs1;r<=grb(2);g<=grb(3);b<=grb(1);

end one;