library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity bigbang is
port(
	clk,rst : in std_logic;
	rxd : in std_logic;
	hs,vs,r,g,b : out std_logic);
end bigbang;

architecture one of bigbang is

signal hs1,vs1,fclk,cclk,sclk : std_logic;
signal fs : std_logic_vector(2 downto 0);
signal cc : std_logic_vector(8 downto 0);
signal ll : std_logic_vector(8 downto 0);
signal grbx : std_logic_vector(3 downto 1);
signal grby : std_logic_vector(3 downto 1);
signal grbp : std_logic_vector(3 downto 1);
signal grb : std_logic_vector(3 downto 1);
signal grbc : std_logic_vector(3 downto 1);
signal mode : std_logic_vector(2 downto 0);

signal clk_cnt,clk_rsclk : std_logic_vector(24 downto 0);
signal PT0,PT1,PT2,PT3,PT4,PT5 : std_logic_vector(3 downto 0);
signal pt : std_logic;

signal freq,scal, sin,tri,squ,rl : std_logic;
type index_type is array(0 to 800) of integer range 0 to 200;
signal tri_ind,squ_ind,sin_ind,sin_id : index_type;
signal x : integer range 0 to 200;
signal sin_y,tri_y,squ_y : integer range 0 to 200;
signal wi : integer range 0 to 7;
signal f,sc : integer range 1 to 8;
signal cci : integer range 0 to 511;
signal rrll : integer range 0 to 200;
signal xt : integer range 0 to 1800;

signal clk_rscnt:integer range 0 to 651;
signal sam_clk:std_logic;
type status_type is(start,data,over);
signal status:status_type;
signal sam_cnt:std_logic_vector(2 downto 0);
signal bit_cnt:std_logic_vector(3 downto 0);
signal rcv_shift_reg:std_logic_vector(7 downto 0);
signal rcv_data:std_logiC_vector(7 downto 0);
signal rrr,l,rot,rev,pul : std_logic;
signal rrrr,uu,lll,dd : std_logic;

type status_stype is array(0 to 17,0 to 17) of std_logic;    --(250-2*2)*(400-4*2)/8=12054--------------64x64--------------
type index_stype is array(0 to 100) of integer range 0 to 127;       --max : 12054--------------4096-------
signal status1,status0 : status_stype;
signal index_x,index_y : index_stype;
signal alive : std_logic;
signal di,dir : std_logic_vector(1 downto 0);
signal i,j,k,m,n : integer range 0 to 127;
signal len : integer range 0 to 100;
signal food : std_logic;
signal food_x,food_y,fx_cnt,fy_cnt : integer range 1 to 16;
signal lcx : std_logic;
signal score1,score0 : std_logic_vector(3 downto 0);
signal ccc,llc : integer range 0 to 127;

type ttstatus_type is array(0 to 11,0 to 42) of std_logic;    --(250-2*2)*(400-4*2)/8=12054
type index_typex is array(0 to 3) of integer range 0 to 15;
type index_typey is array(0 to 3) of integer range 0 to 63;
type tstatuse_type is (start,usual,dead);
signal ttstatus1,ttstatus0 : ttstatus_type;
signal tindex_x : index_typex;
signal tindex_y : index_typey;
signal tstatus : tstatuse_type;
signal food0,food1,food_cnt : integer range 0 to 6;
signal tra,tra_r,tra_l,tra_ro,tra_re,tra_d : std_logic;
signal ti,tj,tk,tm,tn,tsp : integer range 0 to 63;
signal tccc,tlll : integer range 0 to 511;

begin
grb(2)<=(grbp(2))and hs1 and vs1;
grb(3)<=(grbp(3))and hs1 and vs1;
grb(1)<=(grbp(1))and hs1 and vs1;


------------------------------------rs232-------------------------------

P1:process(clk,rst)
begin
	if rst='0' then
		clk_rscnt<=0;
	elsif rising_edge(clk) then
		if clk_rscnt=651 then
			clk_rscnt<=0;
			sam_clk<='1';
		else
			clk_rscnt<=clk_rscnt+1;
			sam_clk<='0';
		end if;
	end if;
end process P1;

P2:process(clk,rst)
begin
	if rst='0' then
		status<=start;
		sam_cnt<="000";
		bit_cnt<="0000";
		rcv_shift_reg<="00111111";
		rcv_data<="00111111";

		freq<='0';
		scal<='0'; 
		sin<='1';
		tri<='1';
		squ<='1';
		rl<='0';
		rrll<=0;

		rrr<='0';
		l<='0';
		rot<='0';
		rev<='0';
		pul<='0';

		rrrr<='0';
		uu<='0';
		lll<='0';
		dd<='0';

	elsif rising_edge(clk) then
		if sam_clk='1' then
			case status is
				when start=>
					if rxd='0' then
						if sam_cnt="011" then
							sam_cnt<="000";
							status<=data;
							bit_cnt<="0000";
						else
							sam_cnt<=sam_cnt+'1';
						end if;
					end if;
				when data=>
					if sam_cnt="111" then
						if bit_cnt="1000" then
							status<=over;
						else
							rcv_shift_reg<=rxd&rcv_shift_reg(7 downto 1);
							sam_cnt<="000";
							bit_cnt<=bit_cnt+'1';
						end if;
					else
						sam_cnt<=sam_cnt+'1';
					end if;
				when over=>
					rcv_data<=rcv_shift_reg;
					
					if rcv_data="00001010" then
						if mode="111" then               
							mode<="000";
						else
							mode<=mode+1;
						end if;		
					end if;	
					mode<="111";	
					if mode="101" then
						if rcv_data="01110001" then
							if f=8 then
							f<=1;
							else
							f<=f+1;
							end if;
						elsif rcv_data="01110111" then
							if sc=8 then
							sc<=1;
							elsif (sc=1 or sc=2 or sc=4) then
							sc<=sc*2;
							else
							sc<=1;
							end if;
						elsif rcv_data="01100101" then
							sin<=not sin;
						elsif rcv_data="01110010" then
							tri<=not tri;
						elsif rcv_data="01110100" then
							squ<=not squ;
						elsif rcv_data="01111001" then
							if rrll=200 then
							rrll<=0;
							else 
							rrll<=rrll+1;
							end if;
						end if;	
						
					elsif mode="111" then
						if rcv_data="01100001" then
							rrr<=not rrr;l<='0';rot<='0';rev<='0';pul<='0';
						elsif rcv_data="01110011" then
							l<=not l;rrr<='0';rot<='0';rev<='0';pul<='0';
						elsif rcv_data="01100100" then
							rot<=not rot;rrr<='0';l<='0';rev<='0';pul<='0';
						elsif rcv_data="01100110" then
							rev<=not rev;rrr<='0';l<='0';rot<='0';pul<='0';
						elsif rcv_data="01100111" then
							pul<=not pul;rrr<='0';l<='0';rot<='0';rev<='0';
						end if;
					elsif mode="110" then
						if rcv_data="01111010" then
							rrrr<=not rrrr;
						elsif rcv_data="01111000" then
							uu<=not uu;
						elsif rcv_data="01100011" then
							lll<=not lll;
						elsif rcv_data="01110110" then
							dd<=not dd;
						end if;
					end if;
					
					status<=start;
			end case;
		end if;
	end if;
end process P2;


    PROCESS( CLK )
    BEGIN
        IF CLK'EVENT AND CLK = '1' THEN -- 50MHz 5分频
            IF FS = 4 THEN FS <= "000";
            ELSE
                FS <= (FS + 1);
            END IF;
        END IF;
    END PROCESS;
    FCLK <= FS(2);
    PROCESS( FCLK )--再315分频，12000000/(13*30)=30769,接近于行频31469
    BEGIN
        IF FCLK'EVENT AND FCLK = '1' THEN
            IF CC = 314 THEN  CC <= "000000000";
            ELSE
                CC <= CC + 1;
            END IF;
        END IF;
    END PROCESS;
    CCLK <= CC(8);
    
    PROCESS( CCLK )
    BEGIN
        IF CCLK'EVENT AND CCLK = '0' THEN
            IF LL = 481 THEN  LL <= "000000000";
            ELSE
                LL <= LL + 1;
            END IF;
        END IF;
    END PROCESS;
    
    
    PROCESS( CC,LL )
    BEGIN
        IF CC > 251 THEN  HS1 <= '0';  --行同步
        ELSE
            HS1 <= '1';
        END IF;
        IF LL > 479 THEN  VS1 <= '0'; --场同步
        ELSE
            VS1 <= '1';
        END IF;
    END PROCESS;
    
process(clk)
begin
	if rising_edge(clk) then
		IF clk_cnt=25000000 THEN clk_cnt<=(others=>'0');
        ELSE
            clk_cnt<=clk_cnt+1;
        END IF;
    END IF;
END PROCESS;

sclk<=clk_cnt(24);
----------------------------------------clk------------------------------
process(sclk,rst)
begin
if rst='0' then

PT0<="0000";PT1<="0000";PT2<="0000";PT3<="0000";PT4<="0000";PT5<="0000";pt<='0';

elsif rising_edge(sclk) then
pt<=not pt;
if pt='1' and pul='0' then
	if PT4="0101" and PT5="1001" then
		if PT2="0101" and PT3="1001" then
			if PT0="0010" and PT1="0011" then
				PT0<="0000";PT1<="0000";
			elsif PT1="1001" then
				PT0<=PT0+1;PT1<="0000";
			else
				PT1<=PT1+1;
			end if;
			PT2<="0000";PT3<="0000";
		elsif PT3="1001" then
			PT2<=PT2+1;PT3<="0000";
		else
			PT3<=PT3+1;
		end if;
		PT4<="0000";PT5<="0000";
	elsif PT5="1001" then
		PT4<=PT4+1;PT5<="0000";
	else
		PT5<=PT5+1;
	end if;
end if;
end if;
end process;

 ------------------------------------------wave---------------------------------   

---------------------snake------------------------

process(clk, rst)
begin

if (rst='0') then

if mode="111" then
	food_cnt<=0;
	for i in 1 to 6 loop
		if clk_cnt(i)='1' then
			food_cnt<=food_cnt+1;
		end if;
	end loop;
	for ti in 0 to 42 loop
		ttstatus1(0,ti)<='1';
		ttstatus0(0,ti)<='1';
		ttstatus1(11,ti)<='1';
		ttstatus0(11,ti)<='1';
	end loop;
	for ti in 1 to 10 loop
		ttstatus1(ti,42)<='1';
		ttstatus0(ti,42)<='1';
	end loop;
	for ti in 1 to 10 loop
		for tj in 0 to 41 loop
			ttstatus1(ti,tj)<='0';
			ttstatus0(ti,tj)<='0';
		end loop;
	end loop;
	for ti in 0 to 3 loop
		tindex_x(ti)<=0;
		tindex_y(ti)<=0;
	end loop;
	tstatus<=start;
end if;	
	
score1<="0000";
score0<="0000";

elsif rising_edge(clk) then

if lcx='0' and sclk='1' then

-------------------------------tetris------------------------
if mode="111" then

case tstatus is
when start=>
	food0<=food_cnt;
	if food_cnt=6 then
		food_cnt<=0;
	else
		food_cnt<=food_cnt+1;
	end  if;
	tra<='0';
	case food1 is
	when 0=>
		tindex_x(0)<=5;
		tindex_y(0)<=1;
		tindex_x(1)<=5;
		tindex_y(1)<=2;
		tindex_x(2)<=5;
		tindex_y(2)<=3;
		tindex_x(3)<=5;
		tindex_y(3)<=4;
		
	when 1=>
		tindex_x(0)<=4;
		tindex_y(0)<=1;
		tindex_x(1)<=4;
		tindex_y(1)<=2;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=6;
		tindex_y(3)<=2;
		
	when 2=>
		tindex_x(0)<=5;
		tindex_y(0)<=1;
		tindex_x(1)<=4;
		tindex_y(1)<=2;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=6;
		tindex_y(3)<=2;
		
	when 3=>
		tindex_x(0)<=6;
		tindex_y(0)<=1;
		tindex_x(1)<=4;
		tindex_y(1)<=2;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=6;
		tindex_y(3)<=2;
		
	when 4=>
		tindex_x(0)<=4;
		tindex_y(0)<=1;
		tindex_x(1)<=5;
		tindex_y(1)<=1;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=6;
		tindex_y(3)<=2;
		
	when 5=>
		tindex_x(0)<=6;
		tindex_y(0)<=1;
		tindex_x(1)<=5;
		tindex_y(1)<=1;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=4;
		tindex_y(3)<=2;
		
	when 6=>
		tindex_x(0)<=5;
		tindex_y(0)<=1;
		tindex_x(1)<=6;
		tindex_y(1)<=1;
		tindex_x(2)<=5;
		tindex_y(2)<=2;
		tindex_x(3)<=6;
		tindex_y(3)<=2;
	
	end case;
	
	tstatus<=usual;

when usual=>
	for ti in 0 to 3 loop
		if ttstatus1(tindex_x(ti),tindex_y(ti))='1' then
			tstatus<=dead;
		end if;
	end loop;
	if food_cnt=6 then
		food_cnt<=0;
	else
		food_cnt<=food_cnt+1;
	end  if;
	if pul='0' then
		tra<='0';
		for ti in 0 to 3 loop
			if ttstatus1(tindex_x(ti),tindex_y(ti)+1)='1' then
				tra<='1';
			end if;
		end loop;
		if tra='0' then
			for ti in 0 to 3 loop
				tindex_y(ti)<=tindex_y(ti)+1;
			end loop;
			for ti in 1 to 10 loop
				for tj in 0 to 41 loop
					if ttstatus1(ti,tj)='0' then
						ttstatus0(ti,tj)<='0';
					end if;
				end loop;
			end loop;
			for ti in 0 to 3 loop
				ttstatus0(tindex_x(ti),tindex_y(ti))<='1';
			end loop;
		else
			for ti in 0 to 3 loop
				ttstatus1(tindex_x(ti),tindex_y(ti)-1)<='1';
				ttstatus0(tindex_x(ti),tindex_y(ti)-1)<='0';
			end loop;
			for ti in 1 to 10 loop
				for tj in 0 to 41 loop
					if ttstatus1(ti,tj)='0' then
						ttstatus0(ti,tj)<='0';
					end if;
				end loop;
			end loop;
	
			for ti in 0 to 3 loop
				for tj in 41 downto 1 loop
					tra_d<='1';
					for tk in 1 to 10 loop
						if ttstatus1(tk,tj)='0' then
							tra_d<='0';
						end if;
					end loop;
					if tra_d='1' then
						for tk in 41 downto 1 loop
							if tk<=tj then
								for tsp in 1 to 10 loop
									ttstatus1(tsp,tk)<=ttstatus1(tsp,tk-1);
								end loop;
							end if;
						end loop;
						if score1="1001" and score0="1001" then
							score1<="0000";
							score0<="0000";
						elsif score0="1001" then
							score1<=score1+1;
							score0<="0000";
						else
							score0<=score0+1;
						end if;
					end if;
				end loop;
			end loop;
			food1<=food0;
			tstatus<=start;
		end if;
	end if;
	
	if tstatus=usual then

		if rrr='1' and pul='0' then
			tra_r<='1';
			for ti in 0 to 3 loop
				if ttstatus1(tindex_x(ti)+2,tindex_y(ti)+1)='1' or ttstatus1(tindex_x(ti)+1,tindex_y(ti)+1)='1' then
					tra_r<='0';
				end if;
			end loop;
			if tra_r='1' then
				for ti in 0 to 3 loop
					tindex_x(ti)<=tindex_x(ti)+1;
				end loop;
				for ti in 1 to 10 loop
					for tj in 0 to 41 loop
						if ttstatus1(ti,tj)='0' then
							ttstatus0(ti,tj)<='0';
						end if;
					end loop;
				end loop;
				for ti in 0 to 3 loop
					ttstatus0(tindex_x(ti),tindex_y(ti))<='1';
				end loop;
			end if;
		end if;

		if l='1' and pul='0' then
			tra_l<='1';
			for ti in 0 to 3 loop
				if ttstatus1(tindex_x(ti)-1,tindex_y(ti)+1)='1' or ttstatus1(tindex_x(ti)-2,tindex_y(ti)+1)='1' then
					tra_l<='0';
				end if;
			end loop;
			if tra_l='1' then
				for ti in 0 to 3 loop
					tindex_x(ti)<=tindex_x(ti)-1;
				end loop;
				for ti in 1 to 10 loop
					for tj in 0 to 41 loop
						if ttstatus1(ti,tj)='0' then
							ttstatus0(ti,tj)<='0';
						end if;
					end loop;
				end loop;
				for ti in 0 to 3 loop
					ttstatus0(tindex_x(ti),tindex_y(ti))<='1';
				end loop;
			end if;
		end if;

		if rot='1' and tra='0' and pul='0' then
			tra_ro<='1';
			for ti in 0 to 3 loop
				if ttstatus1(tindex_x(2)+tindex_y(ti)-tindex_y(2),tindex_y(2)+tindex_x(2)-tindex_x(ti)+2)='1' then
					tra_ro<='0';
				end if;
				if ttstatus1(tindex_x(2)+tindex_x(2)-tindex_x(ti),tindex_y(2)+tindex_y(2)-tindex_y(ti)+2)='1' then
					tra_ro<='0';
				end if;
				if ttstatus1(tindex_x(2)+tindex_y(ti)-tindex_y(2),tindex_y(2)+tindex_x(2)-tindex_x(ti)+1)='1' then
					tra_ro<='0';
				end if;
			end loop;
			if tra_ro='1' then
				for ti in 0 to 3 loop
					if ti/=2 then
						tindex_x(ti)<=tindex_x(2)+tindex_y(ti)-tindex_y(2);
						tindex_y(ti)<=tindex_y(2)+tindex_x(2)-tindex_x(ti)+1;
					end if;
				end loop;
				for ti in 1 to 10 loop
					for tj in 0 to 41 loop
						if ttstatus1(ti,tj)='0' then
							ttstatus0(ti,tj)<='0';
						end if;
					end loop;
				end loop;
				for ti in 0 to 3 loop
					ttstatus0(tindex_x(ti),tindex_y(ti))<='1';
				end loop;
			end if;
		end if;
	
		if rev='1' and tra='0' and pul='0' then
			tra_re<='1';
			for ti in 0 to 3 loop
				if ttstatus1(tindex_x(2)+tindex_y(2)-tindex_y(ti),tindex_y(2)+tindex_x(ti)-tindex_x(2)+1)='1' then
					tra_re<='0';
				end if;
				if ttstatus1(tindex_x(2)+tindex_y(2)-tindex_y(ti),tindex_y(2)+tindex_x(ti)-tindex_x(2)+2)='1' then
					tra_re<='0';
				end if;
				if ttstatus1(tindex_x(2)+tindex_x(2)-tindex_x(ti),tindex_y(2)+tindex_y(2)-tindex_y(ti)+2)='1' then
					tra_re<='0';
				end if;
			end loop;
			
			if tra_re='1' then
				for ti in 0 to 3 loop
					if ti/=2 then
						tindex_x(ti)<=tindex_x(2)+tindex_y(2)-tindex_y(ti);
						tindex_y(ti)<=tindex_y(2)+tindex_x(ti)-tindex_x(2)+1;
					end if;
				end loop;
			
				for ti in 1 to 10 loop
					for tj in 0 to 41 loop
						if ttstatus1(ti,tj)='0' then
							ttstatus0(ti,tj)<='0';
						end if;
					end loop;
				end loop;
				for ti in 0 to 3 loop
					ttstatus0(tindex_x(ti),tindex_y(ti))<='1';
				end loop;
			end if;
		end if;
	end if;
		

when dead=>

end case;
end if;

end if;
lcx<=sclk;	
end if;	

end process;
				
process(cc,ll)
begin 
	grbp<="000";


--------------------------------mode="000"--------------------vertical--------------------

-------------------------------mode="110"--------------------snake---------------------
if mode="110" and alive='1' then
	 if cc>89 and cc<165 and ll>100 and ll<252 then
	 ccc<=to_integer(unsigned(cc-90))/4;
	 llc<=to_integer(unsigned(ll-100))/8;

	if status1(ccc,llc)='1' and status0(ccc,llc)='1' then
		grbp<="010";
	elsif status1(ccc,llc)='0' and status0(ccc,llc)='1' then
		grbp<="101";
	elsif status1(ccc,llc)='1' and status0(ccc,llc)='0' then
		grbp<="011";
	end if;
	 end if;
	----------------------------------snake---------begin----------------------

	if (cc=60 and ll=337) then grbp<="010";
	end if;
	if (ll=337 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=338 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=339 and cc>=38 and cc<40) then grbp<="010";
	end if;
	if (ll=339 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=340 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (ll=340 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=341 and cc>=37 and cc<42) then grbp<="010";
	end if;
	if (ll=341 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=342 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=342 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=343 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=343 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=344 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=344 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=345 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=345 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=346 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (cc=54 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=54 and cc<56) then grbp<="010";
	end if;
	if (ll=346 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=346 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=36 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=347 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=347 and cc>=46 and cc<49) then grbp<="010";
	end if;
	if (ll=347 and cc>=53 and cc<57) then grbp<="010";
	end if;
	if (ll=347 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=347 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=347 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=347) then grbp<="010";
	end if;
	if (cc=36 and ll=348) then grbp<="010";
	end if;
	if (ll=348 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=348 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=348 and cc>=46 and cc<49) then grbp<="010";
	end if;
	if (ll=348 and cc>=52 and cc<57) then grbp<="010";
	end if;
	if (ll=348 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=348 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=348 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=348) then grbp<="010";
	end if;
	if (cc=36 and ll=349) then grbp<="010";
	end if;
	if (ll=349 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=349 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=349 and cc>=46 and cc<50) then grbp<="010";
	end if;
	if (ll=349 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=349 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=349 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=349 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=349) then grbp<="010";
	end if;
	if (cc=36 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=36 and cc<39) then grbp<="010";
	end if;
	if (ll=350 and cc>=43 and cc<50) then grbp<="010";
	end if;
	if (ll=350 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=350 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=350 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=350 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=351 and cc>=36 and cc<39) then grbp<="010";
	end if;
	if (ll=351 and cc>=43 and cc<50) then grbp<="010";
	end if;
	if (ll=351 and cc>=53 and cc<58) then grbp<="010";
	end if;
	if (ll=351 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=351 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=351 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=351) then grbp<="010";
	end if;
	if (ll=351 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=352 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=352 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=352 and cc>=47 and cc<50) then grbp<="010";
	end if;
	if (cc=55 and ll=352) then grbp<="010";
	end if;
	if (ll=352 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=352 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=352 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=352 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=352 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=353 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=353 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=353 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=353 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=353 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=353 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (ll=353 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=353 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=354 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=354 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=354 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=354 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=354 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=354 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (ll=354 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=354 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=355 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (ll=355 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=355 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=355 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=355 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=355 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=355 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=356 and cc>=37 and cc<42) then grbp<="010";
	end if;
	if (ll=356 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=356 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=356 and cc>=53 and cc<58) then grbp<="010";
	end if;
	if (ll=356 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=356 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=357 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (ll=357 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=357 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=357 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=357 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=357 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=358 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (ll=358 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=358 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=358 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=358 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=358 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=358) then grbp<="010";
	end if;
	if (ll=358 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=359 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=359 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=359 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=359 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=359 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=359 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=359) then grbp<="010";
	end if;
	if (ll=359 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=360 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=360 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=360 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=360 and cc>=52 and cc<54) then grbp<="010";
	end if;
	if (ll=360 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=360 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=360 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=360) then grbp<="010";
	end if;
	if (ll=360 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=361 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=361 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=361 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=361 and cc>=52 and cc<54) then grbp<="010";
	end if;
	if (ll=361 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=361 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=361 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=362 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=362 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=362 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=362 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=362 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=362 and cc>=60 and cc<66) then grbp<="010";
	end if;
	if (ll=362 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=363 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=363 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=363 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=363 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=363 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=363 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=363 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=363 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (cc=39 and ll=364) then grbp<="010";
	end if;
	if (ll=364 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=364 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=364 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=364 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=364 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=364 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=364 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=364 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=365 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=365 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=365 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=365 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=365 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=365 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=365 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=365 and cc>=68 and cc<71) then grbp<="010";
	end if;
	if (cc=36 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=366 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=366 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=366 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=366 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=366 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=366 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=367 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=367 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=367 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=367 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=367 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=367 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=367 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=367) then grbp<="010";
	end if;
	if (ll=367 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=368 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=368 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=368 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=368 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=368 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=368 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=368 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=369 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=369 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=369 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=369 and cc>=52 and cc<55) then grbp<="010";
	end if;
	if (ll=369 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=369 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=369 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=369 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=369) then grbp<="010";
	end if;
	if (ll=369 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=370 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=370 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=370 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=370 and cc>=52 and cc<55) then grbp<="010";
	end if;
	if (ll=370 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=370 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=370 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=370 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=370) then grbp<="010";
	end if;
	if (cc=38 and ll=371) then grbp<="010";
	end if;
	if (cc=53 and ll=371) then grbp<="010";
	end if;
	if (cc=70 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=70 and cc<72) then grbp<="010";
	end if;


-------------------------------------snake--------------end-------------------

---------------------------------------time-----------begin-------------------

if cc>123 and cc<127 and ll>341 and ll<348 then
	grbp<="010";
end if;
if cc>123 and cc<127 and ll>362 and ll<369 then
	grbp<="010";
end if;

if PT2="0000" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0001" then
	if (cc>95 and cc<101 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0010" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0011" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0100" then
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0101" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0110" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0111" then
	if (cc>90 and cc<96 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="1000" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="1001" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT3="0000" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0001" then
	if (cc>111 and cc<117 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0010" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0011" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0100" then
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0101" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0110" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0111" then
	if (cc>106 and cc<112 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="1000" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="1001" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT4="0000" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0001" then
	if (cc>133 and cc<139 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0010" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0011" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0100" then
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0101" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0110" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0111" then
	if (cc>128 and cc<134 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="1000" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="1001" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT5="0000" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0001" then
	if (cc>149 and cc<155 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0010" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0011" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0100" then
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0101" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0110" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0111" then
	if (cc>144 and cc<150 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="1000" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="1001" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;



---------------------------------------time-------------end---------------------

--------------------------------------score--------------begin-----------------

if score1="0000" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<188 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>194 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0001" then
	if (cc>188 and cc<194 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0010" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0011" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0100" then
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0101" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0110" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0111" then
	if (cc>183 and cc<189 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="1000" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="1001" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if score0="0000" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<204 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>210 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0001" then
	if (cc>204 and cc<210 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0010" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0011" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0100" then
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0101" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0110" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0111" then
	if (cc>199 and cc<205 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="1000" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="1001" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

--------------------------------------score---------end---------------------------


	---------------------------------------------------------------35-75-90-106-122-128-144-160-183-199-215---------
	---------------------------------------------------------------54-318-335-375--------------------------

end if;

if ((mode="110" and alive='0') or (mode="111" and tstatus=dead)) then

	if (cc=69 and ll=135) then grbp<="010";
	end if;
	if (ll=135 and cc>=69 and cc<71) then grbp<="010";
	end if;
	if (ll=136 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=137 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=138 and cc>=68 and cc<74) then grbp<="010";
	end if;
	if (ll=139 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=140 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=141 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=142 and cc>=66 and cc<74) then grbp<="010";
	end if;
	if (ll=143 and cc>=66 and cc<74) then grbp<="010";
	end if;
	if (ll=144 and cc>=66 and cc<74) then grbp<="010";
	end if;
	if (ll=145 and cc>=66 and cc<74) then grbp<="010";
	end if;
	if (ll=146 and cc>=66 and cc<74) then grbp<="010";
	end if;
	if (ll=147 and cc>=65 and cc<74) then grbp<="010";
	end if;
	if (ll=148 and cc>=65 and cc<74) then grbp<="010";
	end if;
	if (ll=149 and cc>=65 and cc<74) then grbp<="010";
	end if;
	if (ll=150 and cc>=65 and cc<74) then grbp<="010";
	end if;
	if (ll=151 and cc>=65 and cc<74) then grbp<="010";
	end if;
	if (ll=152 and cc>=65 and cc<70) then grbp<="010";
	end if;
	if (ll=152 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=153 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (cc=81 and ll=153) then grbp<="010";
	end if;
	if (ll=153 and cc>=81 and cc<83) then grbp<="010";
	end if;
	if (ll=153 and cc>=93 and cc<95) then grbp<="010";
	end if;
	if (ll=153 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (ll=153 and cc>=109 and cc<111) then grbp<="010";
	end if;
	if (cc=65 and ll=154) then grbp<="010";
	end if;
	if (ll=154 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (ll=154 and cc>=79 and cc<83) then grbp<="010";
	end if;
	if (ll=154 and cc>=93 and cc<95) then grbp<="010";
	end if;
	if (ll=154 and cc>=99 and cc<101) then grbp<="010";
	end if;
	if (ll=154 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=154) then grbp<="010";
	end if;
	if (cc=65 and ll=155) then grbp<="010";
	end if;
	if (ll=155 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (ll=155 and cc>=79 and cc<84) then grbp<="010";
	end if;
	if (ll=155 and cc>=88 and cc<90) then grbp<="010";
	end if;
	if (ll=155 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=155 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=155 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=155) then grbp<="010";
	end if;
	if (cc=65 and ll=156) then grbp<="010";
	end if;
	if (ll=156 and cc>=65 and cc<68) then grbp<="010";
	end if;
	if (ll=156 and cc>=78 and cc<84) then grbp<="010";
	end if;
	if (ll=156 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=156 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=156 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=156 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=156) then grbp<="010";
	end if;
	if (cc=64 and ll=157) then grbp<="010";
	end if;
	if (ll=157 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=157 and cc>=78 and cc<84) then grbp<="010";
	end if;
	if (ll=157 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=157 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=157 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=157 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=157) then grbp<="010";
	end if;
	if (ll=157 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=158 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=158 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=158 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=158 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=158 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=158 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=158) then grbp<="010";
	end if;
	if (ll=158 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=159 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=159 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=159 and cc>=88 and cc<102) then grbp<="010";
	end if;
	if (ll=159 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=159) then grbp<="010";
	end if;
	if (ll=159 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=160 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=160 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=160 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=160 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=160) then grbp<="010";
	end if;
	if (ll=160 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=161 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=161 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=161 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=161 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=161) then grbp<="010";
	end if;
	if (ll=161 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=162 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=162 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=162 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=162 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=162) then grbp<="010";
	end if;
	if (ll=162 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=163 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=163 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=163 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=163 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=163) then grbp<="010";
	end if;
	if (ll=163 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=164 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=164 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=164 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=164 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=164) then grbp<="010";
	end if;
	if (ll=164 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=165 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=165 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=165 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=165 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=165) then grbp<="010";
	end if;
	if (ll=165 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=166 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=166 and cc>=78 and cc<85) then grbp<="010";
	end if;
	if (ll=166 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=166 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=166) then grbp<="010";
	end if;
	if (ll=166 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=167 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=167 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (ll=167 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=167 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=167 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=167 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=168 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=168 and cc>=78 and cc<80) then grbp<="010";
	end if;
	if (ll=168 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=168 and cc>=88 and cc<103) then grbp<="010";
	end if;
	if (ll=168 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=168 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=169 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (cc=82 and ll=169) then grbp<="010";
	end if;
	if (ll=169 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=169 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=169 and cc>=93 and cc<98) then grbp<="010";
	end if;
	if (ll=169 and cc>=99 and cc<103) then grbp<="010";
	end if;
	if (ll=169 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=169 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=170 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (cc=82 and ll=170) then grbp<="010";
	end if;
	if (ll=170 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=170 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=170 and cc>=93 and cc<98) then grbp<="010";
	end if;
	if (ll=170 and cc>=99 and cc<103) then grbp<="010";
	end if;
	if (ll=170 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=170 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=171 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=171 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=171 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=171 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=171 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=171 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=171 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=171 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=172 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=172 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=172 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=172 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=172 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=172 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=172 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=172 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=173 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=173 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=173 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=173 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=173 and cc>=94 and cc<98) then grbp<="010";
	end if;
	if (ll=173 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=173 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=173 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=174 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=174 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=174 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=174 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=174 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=174 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=174 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=174 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=175 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=175 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=175 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=175 and cc>=88 and cc<92) then grbp<="010";
	end if;
	if (ll=175 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=175 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=175 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=175 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=176 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=176 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=176 and cc>=81 and cc<86) then grbp<="010";
	end if;
	if (ll=176 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=176 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=176 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=176 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=176 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=177 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=177 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=177 and cc>=81 and cc<86) then grbp<="010";
	end if;
	if (ll=177 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=177 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=177 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=177 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=177 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=178 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=178 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=178 and cc>=79 and cc<86) then grbp<="010";
	end if;
	if (ll=178 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=178 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=178 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=178 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=178) then grbp<="010";
	end if;
	if (ll=178 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=179 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=179 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=179 and cc>=79 and cc<86) then grbp<="010";
	end if;
	if (ll=179 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=179 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=179 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=179 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=179) then grbp<="010";
	end if;
	if (ll=179 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=180 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=180 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=180 and cc>=78 and cc<86) then grbp<="010";
	end if;
	if (ll=180 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=180 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=180 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=180 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=180) then grbp<="010";
	end if;
	if (ll=180 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=181 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=181 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=181 and cc>=78 and cc<86) then grbp<="010";
	end if;
	if (ll=181 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=181 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=181 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=181 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=181) then grbp<="010";
	end if;
	if (ll=181 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=182 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=182 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=182 and cc>=78 and cc<86) then grbp<="010";
	end if;
	if (ll=182 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=182 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=182 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=182 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=182) then grbp<="010";
	end if;
	if (ll=182 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=183 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=183 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=183 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=183 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=183 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=183 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=183 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=183) then grbp<="010";
	end if;
	if (ll=183 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=184 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=184 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=184 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=184 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=184 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=184 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=184 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=184) then grbp<="010";
	end if;
	if (ll=184 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=185 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=185 and cc>=69 and cc<75) then grbp<="010";
	end if;
	if (ll=185 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=185 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=185 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=185 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=185 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=185) then grbp<="010";
	end if;
	if (ll=185 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=186 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=186 and cc>=70 and cc<75) then grbp<="010";
	end if;
	if (ll=186 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=186 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=186 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=186 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=186 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=187 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=187 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=187 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=187 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=187 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=187 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=187 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=188 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=188 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=188 and cc>=77 and cc<81) then grbp<="010";
	end if;
	if (ll=188 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=188 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=188 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=188 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=188 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=188) then grbp<="010";
	end if;
	if (ll=188 and cc>=111 and cc<115) then grbp<="010";
	end if;
	if (ll=189 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=189 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=189 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=189 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=189 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=189 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=189 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=189 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=189) then grbp<="010";
	end if;
	if (ll=189 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=190 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=190 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=190 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=190 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=190 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=190 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=190 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=190 and cc>=105 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=190) then grbp<="010";
	end if;
	if (ll=190 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=191 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=191 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=191 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=191 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=191 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=191 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=191 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=191 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=192 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=192 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=192 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=192 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=192 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=192 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=192 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=192 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=193 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=193 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=193 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=193 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=193 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=193 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=193 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=193 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=194 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=194 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=194 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=194 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=194 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=194 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=194 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=194 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=195 and cc>=64 and cc<68) then grbp<="010";
	end if;
	if (ll=195 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=195 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=195 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=195 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=195 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=195 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=195 and cc>=105 and cc<108) then grbp<="010";
	end if;
	if (ll=196 and cc>=65 and cc<68) then grbp<="010";
	end if;
	if (ll=196 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=196 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=196 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=196 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=196 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=196 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=196 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=197 and cc>=65 and cc<68) then grbp<="010";
	end if;
	if (ll=197 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=197 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=197 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=197 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=197 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=197 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=197 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=198 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (ll=198 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=198 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=198 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=198 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=198 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=198 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=198 and cc>=105 and cc<109) then grbp<="010";
	end if;
	if (ll=199 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (ll=199 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (ll=199 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=199 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=199 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=199 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=199 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=199 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (ll=200 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=200 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=200 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=200 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=200 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=200 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=200 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (cc=65 and ll=201) then grbp<="010";
	end if;
	if (ll=201 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=201 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=201 and cc>=82 and cc<86) then grbp<="010";
	end if;
	if (ll=201 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=201 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=201 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=201 and cc>=106 and cc<109) then grbp<="010";
	end if;
	if (cc=65 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=202 and cc>=77 and cc<80) then grbp<="010";
	end if;
	if (ll=202 and cc>=81 and cc<86) then grbp<="010";
	end if;
	if (ll=202 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=202 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=202 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=202 and cc>=106 and cc<110) then grbp<="010";
	end if;
	if (ll=202 and cc>=112 and cc<114) then grbp<="010";
	end if;
	if (ll=203 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=203 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=203 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=203 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=203 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=203 and cc>=106 and cc<110) then grbp<="010";
	end if;
	if (ll=203 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=204 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=204 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=204 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=204 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=204 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=204 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=205 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=205 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=205 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=205 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=205 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=205 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=205) then grbp<="010";
	end if;
	if (ll=205 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=206 and cc>=65 and cc<75) then grbp<="010";
	end if;
	if (ll=206 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=206 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=206 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=206 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=206 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=207 and cc>=66 and cc<75) then grbp<="010";
	end if;
	if (ll=207 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=207 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=207 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=207 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=207 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=208 and cc>=66 and cc<75) then grbp<="010";
	end if;
	if (ll=208 and cc>=77 and cc<86) then grbp<="010";
	end if;
	if (ll=208 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=208 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=208 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=208 and cc>=106 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=208) then grbp<="010";
	end if;
	if (ll=208 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=209 and cc>=66 and cc<75) then grbp<="010";
	end if;
	if (ll=209 and cc>=77 and cc<82) then grbp<="010";
	end if;
	if (ll=209 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=209 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=209 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=209 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=209 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=209) then grbp<="010";
	end if;
	if (ll=209 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=210 and cc>=66 and cc<75) then grbp<="010";
	end if;
	if (ll=210 and cc>=77 and cc<82) then grbp<="010";
	end if;
	if (ll=210 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=210 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=210 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=210 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=210 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=211 and cc>=66 and cc<75) then grbp<="010";
	end if;
	if (ll=211 and cc>=77 and cc<82) then grbp<="010";
	end if;
	if (ll=211 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=211 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=211 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=211 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=211 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=212 and cc>=67 and cc<75) then grbp<="010";
	end if;
	if (ll=212 and cc>=77 and cc<82) then grbp<="010";
	end if;
	if (ll=212 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=212 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=212 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=212 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=212 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=213 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=213 and cc>=78 and cc<82) then grbp<="010";
	end if;
	if (ll=213 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=213 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=213 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=213 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=213 and cc>=107 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=111 and cc<114) then grbp<="010";
	end if;
	if (ll=214 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=214 and cc>=78 and cc<82) then grbp<="010";
	end if;
	if (ll=214 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=214 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=214 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=214 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=214 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=215 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=215 and cc>=78 and cc<81) then grbp<="010";
	end if;
	if (ll=215 and cc>=83 and cc<86) then grbp<="010";
	end if;
	if (ll=215 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (ll=215 and cc>=94 and cc<97) then grbp<="010";
	end if;
	if (ll=215 and cc>=100 and cc<103) then grbp<="010";
	end if;
	if (ll=215 and cc>=108 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=215) then grbp<="010";
	end if;
	if (ll=215 and cc>=111 and cc<113) then grbp<="010";
	end if;
	if (ll=216 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (ll=216 and cc>=78 and cc<81) then grbp<="010";
	end if;
	if (ll=216 and cc>=109 and cc<111) then grbp<="010";
	end if;
	if (cc=111 and ll=216) then grbp<="010";
	end if;
	if (cc=69 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=69 and cc<71) then grbp<="010";
	end if;
	if (cc=109 and ll=217) then grbp<="010";
	end if;
	if (ll=217 and cc>=109 and cc<111) then grbp<="010";
	end if;

	if (cc=135 and ll=129) then grbp<="010";
	end if;
	if (ll=129 and cc>=135 and cc<137) then grbp<="010";
	end if;
	if (ll=130 and cc>=135 and cc<138) then grbp<="010";
	end if;
	if (ll=131 and cc>=133 and cc<139) then grbp<="010";
	end if;
	if (ll=131 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=132 and cc>=133 and cc<139) then grbp<="010";
	end if;
	if (ll=132 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=133 and cc>=132 and cc<140) then grbp<="010";
	end if;
	if (ll=133 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=134 and cc>=132 and cc<140) then grbp<="010";
	end if;
	if (ll=134 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=135 and cc>=132 and cc<141) then grbp<="010";
	end if;
	if (ll=135 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=136 and cc>=132 and cc<141) then grbp<="010";
	end if;
	if (ll=136 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=137 and cc>=131 and cc<141) then grbp<="010";
	end if;
	if (ll=137 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=138 and cc>=131 and cc<141) then grbp<="010";
	end if;
	if (ll=138 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=139 and cc>=131 and cc<142) then grbp<="010";
	end if;
	if (ll=139 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=140 and cc>=131 and cc<142) then grbp<="010";
	end if;
	if (ll=140 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=141 and cc>=131 and cc<142) then grbp<="010";
	end if;
	if (ll=141 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=142 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=142 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=143 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=143 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=144 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=144 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=145 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=145 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=146 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=146 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=147 and cc>=130 and cc<143) then grbp<="010";
	end if;
	if (ll=147 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=148 and cc>=130 and cc<135) then grbp<="010";
	end if;
	if (ll=148 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (cc=179 and ll=148) then grbp<="010";
	end if;
	if (cc=182 and ll=148) then grbp<="010";
	end if;
	if (ll=148 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=149 and cc>=130 and cc<135) then grbp<="010";
	end if;
	if (ll=149 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=149 and cc>=163 and cc<166) then grbp<="010";
	end if;
	if (cc=178 and ll=149) then grbp<="010";
	end if;
	if (ll=149 and cc>=178 and cc<180) then grbp<="010";
	end if;
	if (ll=149 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=150 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=150 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=150 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=150 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=150 and cc>=162 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=150) then grbp<="010";
	end if;
	if (cc=173 and ll=150) then grbp<="010";
	end if;
	if (ll=150 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (ll=150 and cc>=178 and cc<181) then grbp<="010";
	end if;
	if (ll=150 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=151 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=151 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=151 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=151 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=151 and cc>=162 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=151) then grbp<="010";
	end if;
	if (cc=173 and ll=151) then grbp<="010";
	end if;
	if (ll=151 and cc>=173 and cc<175) then grbp<="010";
	end if;
	if (ll=151 and cc>=178 and cc<181) then grbp<="010";
	end if;
	if (ll=151 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=152 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=152 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=152 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=152 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=152 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=152) then grbp<="010";
	end if;
	if (ll=152 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=152 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=152 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=152 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=153 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=153 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=153 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=153 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=153 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=153) then grbp<="010";
	end if;
	if (ll=153 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=153 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=153 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=153 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=154 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=154 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=154 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=154 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=154 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=154) then grbp<="010";
	end if;
	if (ll=154 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=154 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=154 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=154 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=155 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=155 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=155 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=155 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=155 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=155) then grbp<="010";
	end if;
	if (ll=155 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=155 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=155 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=155 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=156 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=156 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=156 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=156 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=156 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=156) then grbp<="010";
	end if;
	if (ll=156 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=156 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=156 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=156 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=157 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=157 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=157 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=157 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=157 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=157) then grbp<="010";
	end if;
	if (ll=157 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=157 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=157 and cc>=177 and cc<181) then grbp<="010";
	end if;
	if (ll=157 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=158 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=158 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=158 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=158 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=158 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=158) then grbp<="010";
	end if;
	if (ll=158 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=158 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=158 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=159 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=159 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=159 and cc>=145 and cc<149) then grbp<="010";
	end if;
	if (ll=159 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=159 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=159) then grbp<="010";
	end if;
	if (ll=159 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=159 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=159 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=160 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=160 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=160 and cc>=146 and cc<149) then grbp<="010";
	end if;
	if (ll=160 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=160 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=160) then grbp<="010";
	end if;
	if (ll=160 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=160 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=160 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=161 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=161 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=161 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=161 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=161 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=161) then grbp<="010";
	end if;
	if (ll=161 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=161 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=161 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=162 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=162 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=162 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=162 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=162 and cc>=159 and cc<164) then grbp<="010";
	end if;
	if (ll=162 and cc>=165 and cc<169) then grbp<="010";
	end if;
	if (ll=162 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=162 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=163 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=163 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=163 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=163 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=163 and cc>=159 and cc<164) then grbp<="010";
	end if;
	if (ll=163 and cc>=165 and cc<170) then grbp<="010";
	end if;
	if (ll=163 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=163 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=164 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=164 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=164 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=164 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=164 and cc>=159 and cc<164) then grbp<="010";
	end if;
	if (ll=164 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=164 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=164 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=165 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=165 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=165 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=165 and cc>=153 and cc<157) then grbp<="010";
	end if;
	if (ll=165 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=165 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=165 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=165 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=166 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=166 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=166 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=166 and cc>=153 and cc<156) then grbp<="010";
	end if;
	if (ll=166 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=166 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=166 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=166 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=167 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=167 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=167 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=167 and cc>=153 and cc<156) then grbp<="010";
	end if;
	if (ll=167 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=167 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=167 and cc>=173 and cc<180) then grbp<="010";
	end if;
	if (ll=167 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=168 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=168 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=168 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=168 and cc>=153 and cc<156) then grbp<="010";
	end if;
	if (ll=168 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=168 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=168 and cc>=173 and cc<178) then grbp<="010";
	end if;
	if (ll=168 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=169 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=169 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=169 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=169 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=169 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=169 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=169 and cc>=173 and cc<178) then grbp<="010";
	end if;
	if (ll=169 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=170 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=170 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=170 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=170 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=170 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=170 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=170 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=170 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=171 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=171 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=171 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=171 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=171 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=171 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=171 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=171 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=172 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=172 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=172 and cc>=146 and cc<150) then grbp<="010";
	end if;
	if (ll=172 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=172 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=172 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=172 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=172 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=173 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=173 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=173 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=173 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=173 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=173 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=173 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=173 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=174 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=174 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=174 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=174 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=174 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=174 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=174 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=174 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=175 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=175 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=175 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=175 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=175 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=175) then grbp<="010";
	end if;
	if (ll=175 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=175 and cc>=173 and cc<177) then grbp<="010";
	end if;
	if (ll=175 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=176 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=176 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=176 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=176 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=176 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=176) then grbp<="010";
	end if;
	if (ll=176 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=176 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=176 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=177 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=177 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=177 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=177 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=177 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=177) then grbp<="010";
	end if;
	if (ll=177 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=177 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=177 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=178 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=178 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=178 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=178 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=178 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=178) then grbp<="010";
	end if;
	if (ll=178 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=178 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=178 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=179 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=179 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=179 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=179 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=179 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=179) then grbp<="010";
	end if;
	if (ll=179 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=179 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=179 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=180 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=180 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=180 and cc>=147 and cc<150) then grbp<="010";
	end if;
	if (ll=180 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=180 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=180) then grbp<="010";
	end if;
	if (ll=180 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=180 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=180 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=181 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=181 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=181 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=181 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=181 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=181) then grbp<="010";
	end if;
	if (ll=181 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=181 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=181 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=182 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=182 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=182 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=182 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=182 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=182) then grbp<="010";
	end if;
	if (ll=182 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=182 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=182 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=183 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=183 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=183 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=183 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=183 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=183) then grbp<="010";
	end if;
	if (ll=183 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=183 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=183 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=184 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=184 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=184 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=184 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=184 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=184) then grbp<="010";
	end if;
	if (ll=184 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=184 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=184 and cc>=182 and cc<185) then grbp<="010";
	end if;
	if (ll=185 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=185 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=185 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=185 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=185 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=185) then grbp<="010";
	end if;
	if (ll=185 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=185 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=186 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=186 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=186 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=186 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=186 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=186) then grbp<="010";
	end if;
	if (ll=186 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=186 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=187 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=187 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=187 and cc>=147 and cc<151) then grbp<="010";
	end if;
	if (ll=187 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=187 and cc>=159 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=187) then grbp<="010";
	end if;
	if (ll=187 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=187 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=188 and cc>=129 and cc<133) then grbp<="010";
	end if;
	if (ll=188 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=188 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=188 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=188 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=189 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=189 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=189 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=189 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=189 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=190 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=190 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=190 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=190 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=190 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=191 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=191 and cc>=139 and cc<143) then grbp<="010";
	end if;
	if (ll=191 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=191 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=191 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=192 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=192 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=192 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=192 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=192 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=193 and cc>=129 and cc<134) then grbp<="010";
	end if;
	if (ll=193 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=193 and cc>=148 and cc<155) then grbp<="010";
	end if;
	if (ll=193 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=193 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=194 and cc>=130 and cc<134) then grbp<="010";
	end if;
	if (ll=194 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=194 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=194 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=194 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=195 and cc>=130 and cc<135) then grbp<="010";
	end if;
	if (ll=195 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=195 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=195 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=195 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=195 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (ll=196 and cc>=130 and cc<135) then grbp<="010";
	end if;
	if (ll=196 and cc>=138 and cc<143) then grbp<="010";
	end if;
	if (ll=196 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=196 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (ll=196 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=196 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (ll=197 and cc>=130 and cc<143) then grbp<="010";
	end if;
	if (ll=197 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=197 and cc>=159 and cc<163) then grbp<="010";
	end if;
	if (cc=173 and ll=197) then grbp<="010";
	end if;
	if (ll=197 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=197 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=198 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=198 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=198 and cc>=159 and cc<164) then grbp<="010";
	end if;
	if (cc=173 and ll=198) then grbp<="010";
	end if;
	if (ll=198 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=198 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=199 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=199 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=199 and cc>=159 and cc<164) then grbp<="010";
	end if;
	if (ll=199 and cc>=167 and cc<169) then grbp<="010";
	end if;
	if (ll=199 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=199 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=200 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=200 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=200 and cc>=159 and cc<165) then grbp<="010";
	end if;
	if (ll=200 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=200 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=200 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=201 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=201 and cc>=148 and cc<154) then grbp<="010";
	end if;
	if (ll=201 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=201) then grbp<="010";
	end if;
	if (ll=201 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=201 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=201 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=202 and cc>=130 and cc<142) then grbp<="010";
	end if;
	if (ll=202 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=202 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=202) then grbp<="010";
	end if;
	if (ll=202 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=202 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=202 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=203 and cc>=131 and cc<142) then grbp<="010";
	end if;
	if (ll=203 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=203 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=203) then grbp<="010";
	end if;
	if (ll=203 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=203 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=203 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=204 and cc>=131 and cc<142) then grbp<="010";
	end if;
	if (ll=204 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=204 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=204) then grbp<="010";
	end if;
	if (ll=204 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=204 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=204 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=205 and cc>=131 and cc<141) then grbp<="010";
	end if;
	if (ll=205 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=205 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=205) then grbp<="010";
	end if;
	if (ll=205 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=205 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=205 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=206 and cc>=131 and cc<141) then grbp<="010";
	end if;
	if (ll=206 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=206 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=206) then grbp<="010";
	end if;
	if (ll=206 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=206 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=206 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=207 and cc>=131 and cc<141) then grbp<="010";
	end if;
	if (ll=207 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=207 and cc>=160 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=207) then grbp<="010";
	end if;
	if (ll=207 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=207 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=207 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=208 and cc>=132 and cc<141) then grbp<="010";
	end if;
	if (ll=208 and cc>=149 and cc<154) then grbp<="010";
	end if;
	if (ll=208 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=208) then grbp<="010";
	end if;
	if (ll=208 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=208 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=208 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=209 and cc>=132 and cc<141) then grbp<="010";
	end if;
	if (ll=209 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=209 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=209) then grbp<="010";
	end if;
	if (ll=209 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=209 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=209 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=210 and cc>=132 and cc<140) then grbp<="010";
	end if;
	if (ll=210 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=210 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=210) then grbp<="010";
	end if;
	if (ll=210 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=210 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=210 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=211 and cc>=133 and cc<140) then grbp<="010";
	end if;
	if (ll=211 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=211 and cc>=161 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=211) then grbp<="010";
	end if;
	if (ll=211 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=211 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=211 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=212 and cc>=133 and cc<139) then grbp<="010";
	end if;
	if (ll=212 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=212 and cc>=162 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=212) then grbp<="010";
	end if;
	if (ll=212 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=212 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=212 and cc>=182 and cc<186) then grbp<="010";
	end if;
	if (ll=213 and cc>=133 and cc<139) then grbp<="010";
	end if;
	if (ll=213 and cc>=149 and cc<153) then grbp<="010";
	end if;
	if (ll=213 and cc>=162 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=213) then grbp<="010";
	end if;
	if (ll=213 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=213 and cc>=173 and cc<176) then grbp<="010";
	end if;
	if (ll=213 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (ll=214 and cc>=135 and cc<138) then grbp<="010";
	end if;
	if (ll=214 and cc>=163 and cc<166) then grbp<="010";
	end if;
	if (cc=166 and ll=214) then grbp<="010";
	end if;
	if (cc=183 and ll=214) then grbp<="010";
	end if;
	if (ll=214 and cc>=183 and cc<185) then grbp<="010";
	end if;
	if (ll=215 and cc>=135 and cc<137) then grbp<="010";
	end if;
	if (ll=215 and cc>=164 and cc<166) then grbp<="010";
	end if;

	if (cc=65 and ll=230) then grbp<="010";
	end if;
	if (ll=230 and cc>=65 and cc<68) then grbp<="010";
	end if;
	if (ll=230 and cc>=72 and cc<76) then grbp<="010";
	end if;
	if (ll=231 and cc>=65 and cc<69) then grbp<="010";
	end if;
	if (ll=231 and cc>=72 and cc<76) then grbp<="010";
	end if;
	if (ll=232 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=232 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=233 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=233 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=234 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=234 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=235 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=235 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=236 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=236 and cc>=72 and cc<75) then grbp<="010";
	end if;
	if (ll=237 and cc>=66 and cc<69) then grbp<="010";
	end if;
	if (ll=237 and cc>=71 and cc<75) then grbp<="010";
	end if;
	if (cc=103 and ll=237) then grbp<="010";
	end if;
	if (cc=66 and ll=238) then grbp<="010";
	end if;
	if (ll=238 and cc>=66 and cc<70) then grbp<="010";
	end if;
	if (ll=238 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=238 and cc>=78 and cc<82) then grbp<="010";
	end if;
	if (ll=238 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=238 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=238 and cc>=98 and cc<100) then grbp<="010";
	end if;
	if (ll=238 and cc>=102 and cc<104) then grbp<="010";
	end if;
	if (ll=239 and cc>=67 and cc<70) then grbp<="010";
	end if;
	if (ll=239 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=239 and cc>=78 and cc<83) then grbp<="010";
	end if;
	if (ll=239 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=239 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=239 and cc>=98 and cc<100) then grbp<="010";
	end if;
	if (ll=239 and cc>=102 and cc<104) then grbp<="010";
	end if;
	if (ll=240 and cc>=67 and cc<70) then grbp<="010";
	end if;
	if (ll=240 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=240 and cc>=77 and cc<83) then grbp<="010";
	end if;
	if (ll=240 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=240 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=240 and cc>=98 and cc<100) then grbp<="010";
	end if;
	if (ll=240 and cc>=101 and cc<104) then grbp<="010";
	end if;
	if (ll=241 and cc>=67 and cc<70) then grbp<="010";
	end if;
	if (ll=241 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=241 and cc>=77 and cc<84) then grbp<="010";
	end if;
	if (ll=241 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=241 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=241 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=242 and cc>=67 and cc<70) then grbp<="010";
	end if;
	if (ll=242 and cc>=71 and cc<74) then grbp<="010";
	end if;
	if (ll=242 and cc>=77 and cc<84) then grbp<="010";
	end if;
	if (ll=242 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=242 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=242 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=243 and cc>=67 and cc<74) then grbp<="010";
	end if;
	if (ll=243 and cc>=76 and cc<84) then grbp<="010";
	end if;
	if (ll=243 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=243 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=243 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=244 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=244 and cc>=76 and cc<84) then grbp<="010";
	end if;
	if (ll=244 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=244 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=244 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=245 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=245 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=245 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (ll=245 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=245 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=245 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=246 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=246 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=246 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (ll=246 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=246 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=246 and cc>=98 and cc<104) then grbp<="010";
	end if;
	if (ll=247 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=247 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=247 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (ll=247 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=247 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=247 and cc>=98 and cc<102) then grbp<="010";
	end if;
	if (ll=248 and cc>=68 and cc<73) then grbp<="010";
	end if;
	if (ll=248 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=248 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=248 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=248 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=248 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=249 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (ll=249 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=249 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=249 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=249 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=249 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=250 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (ll=250 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=250 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=250 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=250 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=250 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=251 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=251 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=251 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=251 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=251 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=251 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=252 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=252 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=252 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=252 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=252 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=252 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=253 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=253 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=253 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=253 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=253 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=253 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=254 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=254 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=254 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=254 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=254 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=254 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=255 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=255 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=255 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=255 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=255 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=255 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=256 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=256 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=256 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=256 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=256 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=256 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=257 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=257 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=257 and cc>=82 and cc<85) then grbp<="010";
	end if;
	if (ll=257 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=257 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=257 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=258 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=258 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=258 and cc>=81 and cc<85) then grbp<="010";
	end if;
	if (ll=258 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=258 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=258 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=259 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=259 and cc>=76 and cc<79) then grbp<="010";
	end if;
	if (ll=259 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (ll=259 and cc>=87 and cc<90) then grbp<="010";
	end if;
	if (ll=259 and cc>=92 and cc<96) then grbp<="010";
	end if;
	if (ll=259 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=260 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=260 and cc>=76 and cc<80) then grbp<="010";
	end if;
	if (ll=260 and cc>=81 and cc<84) then grbp<="010";
	end if;
	if (ll=260 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (ll=260 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=261 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=261 and cc>=76 and cc<84) then grbp<="010";
	end if;
	if (ll=261 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (ll=261 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=262 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=262 and cc>=77 and cc<84) then grbp<="010";
	end if;
	if (ll=262 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (ll=262 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=263 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=263 and cc>=77 and cc<84) then grbp<="010";
	end if;
	if (ll=263 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (ll=263 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=264 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=264 and cc>=77 and cc<83) then grbp<="010";
	end if;
	if (ll=264 and cc>=87 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=91 and cc<96) then grbp<="010";
	end if;
	if (ll=264 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=265 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=265 and cc>=78 and cc<83) then grbp<="010";
	end if;
	if (ll=265 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=265) then grbp<="010";
	end if;
	if (cc=93 and ll=265) then grbp<="010";
	end if;
	if (ll=265 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=265 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=266 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (ll=266 and cc>=78 and cc<82) then grbp<="010";
	end if;
	if (ll=266 and cc>=88 and cc<91) then grbp<="010";
	end if;
	if (cc=91 and ll=266) then grbp<="010";
	end if;
	if (cc=93 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=93 and cc<96) then grbp<="010";
	end if;
	if (ll=266 and cc>=98 and cc<101) then grbp<="010";
	end if;
	if (ll=267 and cc>=79 and cc<81) then grbp<="010";
	end if;
	if (ll=267 and cc>=89 and cc<91) then grbp<="010";
	end if;






	if (cc=65 and ll=229) then grbp<="111";
	end if;
	if (ll=229 and cc>=65 and cc<105) then grbp<="111";
	end if;
	if (cc=68 and ll=230) then grbp<="111";
	end if;
	if (ll=230 and cc>=68 and cc<72) then grbp<="111";
	end if;
	if (ll=230 and cc>=76 and cc<105) then grbp<="111";
	end if;
	if (cc=69 and ll=231) then grbp<="111";
	end if;
	if (ll=231 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=231 and cc>=76 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=232) then grbp<="111";
	end if;
	if (cc=69 and ll=232) then grbp<="111";
	end if;
	if (ll=232 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=232 and cc>=75 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=233) then grbp<="111";
	end if;
	if (cc=69 and ll=233) then grbp<="111";
	end if;
	if (ll=233 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=233 and cc>=75 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=234) then grbp<="111";
	end if;
	if (cc=69 and ll=234) then grbp<="111";
	end if;
	if (ll=234 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=234 and cc>=75 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=235) then grbp<="111";
	end if;
	if (cc=69 and ll=235) then grbp<="111";
	end if;
	if (ll=235 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=235 and cc>=75 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=236) then grbp<="111";
	end if;
	if (cc=69 and ll=236) then grbp<="111";
	end if;
	if (ll=236 and cc>=69 and cc<72) then grbp<="111";
	end if;
	if (ll=236 and cc>=75 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=237) then grbp<="111";
	end if;
	if (cc=69 and ll=237) then grbp<="111";
	end if;
	if (ll=237 and cc>=69 and cc<71) then grbp<="111";
	end if;
	if (ll=237 and cc>=75 and cc<80) then grbp<="111";
	end if;
	if (ll=237 and cc>=81 and cc<103) then grbp<="111";
	end if;
	if (cc=65 and ll=238) then grbp<="111";
	end if;
	if (cc=70 and ll=238) then grbp<="111";
	end if;
	if (cc=74 and ll=238) then grbp<="111";
	end if;
	if (ll=238 and cc>=74 and cc<78) then grbp<="111";
	end if;
	if (ll=238 and cc>=82 and cc<87) then grbp<="111";
	end if;
	if (ll=238 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=238 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=238 and cc>=100 and cc<102) then grbp<="111";
	end if;
	if (cc=65 and ll=239) then grbp<="111";
	end if;
	if (ll=239 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (cc=74 and ll=239) then grbp<="111";
	end if;
	if (ll=239 and cc>=74 and cc<78) then grbp<="111";
	end if;
	if (ll=239 and cc>=83 and cc<87) then grbp<="111";
	end if;
	if (ll=239 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=239 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=239 and cc>=100 and cc<102) then grbp<="111";
	end if;
	if (cc=65 and ll=240) then grbp<="111";
	end if;
	if (ll=240 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (cc=74 and ll=240) then grbp<="111";
	end if;
	if (ll=240 and cc>=74 and cc<77) then grbp<="111";
	end if;
	if (ll=240 and cc>=83 and cc<87) then grbp<="111";
	end if;
	if (ll=240 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=240 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=104 and ll=240) then grbp<="111";
	end if;
	if (cc=65 and ll=241) then grbp<="111";
	end if;
	if (ll=241 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (cc=74 and ll=241) then grbp<="111";
	end if;
	if (ll=241 and cc>=74 and cc<77) then grbp<="111";
	end if;
	if (ll=241 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=241 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=241 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=242) then grbp<="111";
	end if;
	if (ll=242 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (cc=74 and ll=242) then grbp<="111";
	end if;
	if (ll=242 and cc>=74 and cc<77) then grbp<="111";
	end if;
	if (ll=242 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=242 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=242 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=243) then grbp<="111";
	end if;
	if (ll=243 and cc>=65 and cc<67) then grbp<="111";
	end if;
	if (ll=243 and cc>=74 and cc<76) then grbp<="111";
	end if;
	if (ll=243 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=243 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=243 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=244) then grbp<="111";
	end if;
	if (ll=244 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=244 and cc>=73 and cc<76) then grbp<="111";
	end if;
	if (ll=244 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=244 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=244 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=245) then grbp<="111";
	end if;
	if (ll=245 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=245 and cc>=73 and cc<76) then grbp<="111";
	end if;
	if (ll=245 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=245 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=245 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=245 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=246) then grbp<="111";
	end if;
	if (ll=246 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=246 and cc>=73 and cc<76) then grbp<="111";
	end if;
	if (ll=246 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=246 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=246 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=246 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (cc=65 and ll=247) then grbp<="111";
	end if;
	if (ll=247 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=247 and cc>=73 and cc<76) then grbp<="111";
	end if;
	if (ll=247 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=247 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=247 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=247 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=247 and cc>=102 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=248) then grbp<="111";
	end if;
	if (ll=248 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=248 and cc>=73 and cc<76) then grbp<="111";
	end if;
	if (ll=248 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=248 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=248 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=248 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=248 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=249) then grbp<="111";
	end if;
	if (ll=249 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=249 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=249 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=249 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=249 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=249 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=249 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=250) then grbp<="111";
	end if;
	if (ll=250 and cc>=65 and cc<68) then grbp<="111";
	end if;
	if (ll=250 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=250 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=250 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=250 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=250 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=250 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=251) then grbp<="111";
	end if;
	if (ll=251 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=251 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=251 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=251 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=251 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=251 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=251 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=252) then grbp<="111";
	end if;
	if (ll=252 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=252 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=252 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=252 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=252 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=252 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=252 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=253) then grbp<="111";
	end if;
	if (ll=253 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=253 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=253 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=253 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=253 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=253 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=253 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=254) then grbp<="111";
	end if;
	if (ll=254 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=254 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=254 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=254 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=254 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=254 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=254 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=255) then grbp<="111";
	end if;
	if (ll=255 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=255 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=255 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=255 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=255 and cc>=90 and cc<93) then grbp<="111";
	end if;
	if (ll=255 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=255 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=256) then grbp<="111";
	end if;
	if (ll=256 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=256 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=256 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=256 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=256 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (ll=256 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=256 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=257) then grbp<="111";
	end if;
	if (ll=257 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=257 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=257 and cc>=79 and cc<82) then grbp<="111";
	end if;
	if (ll=257 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=257 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (ll=257 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=257 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=258) then grbp<="111";
	end if;
	if (ll=258 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=258 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=258 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=258 and cc>=85 and cc<87) then grbp<="111";
	end if;
	if (ll=258 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (ll=258 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=258 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=259) then grbp<="111";
	end if;
	if (ll=259 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=259 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=259 and cc>=79 and cc<81) then grbp<="111";
	end if;
	if (ll=259 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=259 and cc>=90 and cc<92) then grbp<="111";
	end if;
	if (ll=259 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=259 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=260 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (cc=84 and ll=260) then grbp<="111";
	end if;
	if (ll=260 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=260 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=260 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=261) then grbp<="111";
	end if;
	if (ll=261 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=261 and cc>=72 and cc<76) then grbp<="111";
	end if;
	if (ll=261 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=261 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=261 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=262) then grbp<="111";
	end if;
	if (ll=262 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=262 and cc>=72 and cc<77) then grbp<="111";
	end if;
	if (ll=262 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=262 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=262 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=263) then grbp<="111";
	end if;
	if (ll=263 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=263 and cc>=72 and cc<77) then grbp<="111";
	end if;
	if (ll=263 and cc>=84 and cc<87) then grbp<="111";
	end if;
	if (ll=263 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=263 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=264) then grbp<="111";
	end if;
	if (ll=264 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=264 and cc>=72 and cc<77) then grbp<="111";
	end if;
	if (ll=264 and cc>=83 and cc<87) then grbp<="111";
	end if;
	if (ll=264 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=264 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=265 and cc>=72 and cc<78) then grbp<="111";
	end if;
	if (ll=265 and cc>=83 and cc<88) then grbp<="111";
	end if;
	if (cc=96 and ll=265) then grbp<="111";
	end if;
	if (ll=265 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=265 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=266) then grbp<="111";
	end if;
	if (ll=266 and cc>=65 and cc<69) then grbp<="111";
	end if;
	if (ll=266 and cc>=72 and cc<78) then grbp<="111";
	end if;
	if (ll=266 and cc>=82 and cc<88) then grbp<="111";
	end if;
	if (cc=96 and ll=266) then grbp<="111";
	end if;
	if (ll=266 and cc>=96 and cc<98) then grbp<="111";
	end if;
	if (ll=266 and cc>=101 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=267) then grbp<="111";
	end if;
	if (ll=267 and cc>=65 and cc<79) then grbp<="111";
	end if;
	if (ll=267 and cc>=81 and cc<89) then grbp<="111";
	end if;
	if (ll=267 and cc>=91 and cc<105) then grbp<="111";
	end if;
	if (cc=65 and ll=268) then grbp<="111";
	end if;
	if (ll=268 and cc>=65 and cc<105) then grbp<="111";
	end if;

	if (cc=117 and ll=229) then grbp<="010";
	end if;
	if (ll=229 and cc>=117 and cc<120) then grbp<="010";
	end if;
	if (ll=230 and cc>=116 and cc<121) then grbp<="010";
	end if;
	if (ll=231 and cc>=115 and cc<122) then grbp<="010";
	end if;
	if (ll=232 and cc>=115 and cc<122) then grbp<="010";
	end if;
	if (ll=233 and cc>=115 and cc<122) then grbp<="010";
	end if;
	if (ll=234 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=235 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=236 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=237 and cc>=114 and cc<118) then grbp<="010";
	end if;
	if (ll=237 and cc>=119 and cc<121) then grbp<="010";
	end if;
	if (ll=238 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (cc=127 and ll=238) then grbp<="010";
	end if;
	if (ll=238 and cc>=127 and cc<130) then grbp<="010";
	end if;
	if (ll=238 and cc>=136 and cc<139) then grbp<="010";
	end if;
	if (ll=238 and cc>=144 and cc<146) then grbp<="010";
	end if;
	if (ll=238 and cc>=149 and cc<151) then grbp<="010";
	end if;
	if (ll=238 and cc>=154 and cc<158) then grbp<="010";
	end if;
	if (cc=114 and ll=239) then grbp<="010";
	end if;
	if (ll=239 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (ll=239 and cc>=126 and cc<131) then grbp<="010";
	end if;
	if (ll=239 and cc>=135 and cc<140) then grbp<="010";
	end if;
	if (ll=239 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=239 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=239 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=239) then grbp<="010";
	end if;
	if (cc=114 and ll=240) then grbp<="010";
	end if;
	if (ll=240 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (ll=240 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=240 and cc>=134 and cc<140) then grbp<="010";
	end if;
	if (ll=240 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=240 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=240 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=240) then grbp<="010";
	end if;
	if (cc=114 and ll=241) then grbp<="010";
	end if;
	if (ll=241 and cc>=114 and cc<117) then grbp<="010";
	end if;
	if (ll=241 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=241 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=241 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=241 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=241 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=241) then grbp<="010";
	end if;
	if (cc=114 and ll=242) then grbp<="010";
	end if;
	if (ll=242 and cc>=114 and cc<118) then grbp<="010";
	end if;
	if (ll=242 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=242 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=242 and cc>=144 and cc<151) then grbp<="010";
	end if;
	if (ll=242 and cc>=152 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=242) then grbp<="010";
	end if;
	if (ll=242 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=243 and cc>=114 and cc<118) then grbp<="010";
	end if;
	if (ll=243 and cc>=124 and cc<131) then grbp<="010";
	end if;
	if (ll=243 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=243 and cc>=144 and cc<150) then grbp<="010";
	end if;
	if (ll=243 and cc>=152 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=243) then grbp<="010";
	end if;
	if (ll=243 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=244 and cc>=114 and cc<119) then grbp<="010";
	end if;
	if (ll=244 and cc>=124 and cc<131) then grbp<="010";
	end if;
	if (ll=244 and cc>=133 and cc<141) then grbp<="010";
	end if;
	if (ll=244 and cc>=144 and cc<150) then grbp<="010";
	end if;
	if (ll=244 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=244 and cc>=157 and cc<160) then grbp<="010";
	end if;
	if (ll=245 and cc>=114 and cc<119) then grbp<="010";
	end if;
	if (ll=245 and cc>=124 and cc<128) then grbp<="010";
	end if;
	if (ll=245 and cc>=129 and cc<131) then grbp<="010";
	end if;
	if (ll=245 and cc>=133 and cc<137) then grbp<="010";
	end if;
	if (ll=245 and cc>=138 and cc<142) then grbp<="010";
	end if;
	if (ll=245 and cc>=144 and cc<150) then grbp<="010";
	end if;
	if (ll=245 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=245 and cc>=157 and cc<160) then grbp<="010";
	end if;
	if (ll=246 and cc>=114 and cc<120) then grbp<="010";
	end if;
	if (ll=246 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (cc=133 and ll=246) then grbp<="010";
	end if;
	if (ll=246 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=246 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=246 and cc>=144 and cc<150) then grbp<="010";
	end if;
	if (ll=246 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=246 and cc>=157 and cc<160) then grbp<="010";
	end if;
	if (ll=247 and cc>=115 and cc<121) then grbp<="010";
	end if;
	if (ll=247 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=247 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=247 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=247 and cc>=144 and cc<148) then grbp<="010";
	end if;
	if (ll=247 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=247 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=248 and cc>=115 and cc<121) then grbp<="010";
	end if;
	if (ll=248 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=248 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=248 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=248 and cc>=144 and cc<148) then grbp<="010";
	end if;
	if (ll=248 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=248 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=249 and cc>=115 and cc<121) then grbp<="010";
	end if;
	if (ll=249 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=249 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=249 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=249 and cc>=144 and cc<148) then grbp<="010";
	end if;
	if (ll=249 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=249 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=250 and cc>=116 and cc<122) then grbp<="010";
	end if;
	if (ll=250 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=250 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=250 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=250 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=250 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=250) then grbp<="010";
	end if;
	if (ll=250 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=251 and cc>=116 and cc<122) then grbp<="010";
	end if;
	if (ll=251 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=251 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=251 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=251 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=251 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=251) then grbp<="010";
	end if;
	if (ll=251 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=252 and cc>=117 and cc<122) then grbp<="010";
	end if;
	if (ll=252 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=252 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=252 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=252 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=252 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=252) then grbp<="010";
	end if;
	if (ll=252 and cc>=158 and cc<161) then grbp<="010";
	end if;
	if (ll=253 and cc>=118 and cc<122) then grbp<="010";
	end if;
	if (ll=253 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=253 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=253 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=253 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=253 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=253) then grbp<="010";
	end if;
	if (ll=253 and cc>=158 and cc<161) then grbp<="010";
	end if;
	if (ll=254 and cc>=118 and cc<122) then grbp<="010";
	end if;
	if (ll=254 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=254 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=254 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=254 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=254 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=254) then grbp<="010";
	end if;
	if (ll=254 and cc>=158 and cc<161) then grbp<="010";
	end if;
	if (ll=255 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (ll=255 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=255 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=255 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=255 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=255 and cc>=151 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=255) then grbp<="010";
	end if;
	if (ll=255 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=256 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (ll=256 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=256 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=256 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=256 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=256 and cc>=151 and cc<155) then grbp<="010";
	end if;
	if (ll=257 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (ll=257 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=257 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=257 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=257 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=257 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=258 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (ll=258 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=258 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=258 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=258 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=258 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (cc=119 and ll=259) then grbp<="010";
	end if;
	if (ll=259 and cc>=119 and cc<122) then grbp<="010";
	end if;
	if (ll=259 and cc>=124 and cc<127) then grbp<="010";
	end if;
	if (ll=259 and cc>=133 and cc<136) then grbp<="010";
	end if;
	if (ll=259 and cc>=139 and cc<142) then grbp<="010";
	end if;
	if (ll=259 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=259 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (ll=260 and cc>=114 and cc<116) then grbp<="010";
	end if;
	if (ll=260 and cc>=118 and cc<122) then grbp<="010";
	end if;
	if (ll=260 and cc>=124 and cc<128) then grbp<="010";
	end if;
	if (cc=133 and ll=260) then grbp<="010";
	end if;
	if (ll=260 and cc>=133 and cc<137) then grbp<="010";
	end if;
	if (ll=260 and cc>=138 and cc<142) then grbp<="010";
	end if;
	if (ll=260 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=260 and cc>=152 and cc<155) then grbp<="010";
	end if;
	if (cc=114 and ll=261) then grbp<="010";
	end if;
	if (ll=261 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=261 and cc>=124 and cc<131) then grbp<="010";
	end if;
	if (ll=261 and cc>=133 and cc<142) then grbp<="010";
	end if;
	if (ll=261 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=261 and cc>=152 and cc<156) then grbp<="010";
	end if;
	if (ll=261 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=262 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=262 and cc>=124 and cc<131) then grbp<="010";
	end if;
	if (ll=262 and cc>=133 and cc<141) then grbp<="010";
	end if;
	if (ll=262 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=262 and cc>=152 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=262) then grbp<="010";
	end if;
	if (ll=262 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=263 and cc>=114 and cc<122) then grbp<="010";
	end if;
	if (ll=263 and cc>=124 and cc<131) then grbp<="010";
	end if;
	if (ll=263 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=263 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=263 and cc>=152 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=263) then grbp<="010";
	end if;
	if (ll=263 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=264 and cc>=114 and cc<121) then grbp<="010";
	end if;
	if (ll=264 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=264 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=264 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=264 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=264) then grbp<="010";
	end if;
	if (ll=264 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=265 and cc>=114 and cc<121) then grbp<="010";
	end if;
	if (ll=265 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=265 and cc>=134 and cc<141) then grbp<="010";
	end if;
	if (ll=265 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=265 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=265) then grbp<="010";
	end if;
	if (ll=265 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=266 and cc>=114 and cc<120) then grbp<="010";
	end if;
	if (ll=266 and cc>=125 and cc<131) then grbp<="010";
	end if;
	if (ll=266 and cc>=135 and cc<140) then grbp<="010";
	end if;
	if (ll=266 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=266 and cc>=153 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=266) then grbp<="010";
	end if;
	if (ll=266 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=267 and cc>=115 and cc<120) then grbp<="010";
	end if;
	if (ll=267 and cc>=126 and cc<130) then grbp<="010";
	end if;
	if (ll=267 and cc>=135 and cc<140) then grbp<="010";
	end if;
	if (ll=267 and cc>=144 and cc<147) then grbp<="010";
	end if;
	if (ll=267 and cc>=154 and cc<158) then grbp<="010";
	end if;
	if (cc=158 and ll=267) then grbp<="010";
	end if;
	if (cc=116 and ll=268) then grbp<="010";
	end if;
	if (ll=268 and cc>=116 and cc<119) then grbp<="010";
	end if;
	if (ll=268 and cc>=127 and cc<129) then grbp<="010";
	end if;
	if (ll=268 and cc>=136 and cc<139) then grbp<="010";
	end if;
	if (ll=268 and cc>=155 and cc<158) then grbp<="010";
	end if;

if score1="0000" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>169 and cc<172 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>175 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0001" then
	if (cc>172 and cc<175 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0010" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0011" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0100" then
	if (cc>169 and cc<173 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0101" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0110" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="0111" then
	if (cc>169 and cc<173 and ll>227 and ll<232) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score1="1000" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score1="1001" then
	if (cc>169 and cc<178 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>169 and cc<173 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>174 and cc<178 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>169 and cc<178 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;

if score0="0000" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>178 and cc<181 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>184 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0001" then
	if (cc>181 and cc<184 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0010" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<182 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0011" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0100" then
	if (cc>178 and cc<182 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0101" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>178 and cc<182 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0110" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>178 and cc<182 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>245 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="0111" then
	if (cc>178 and cc<182 and ll>227 and ll<232) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
end if;
if score0="1000" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>178 and cc<182 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;
if score0="1001" then
	if (cc>178 and cc<187 and ll>227 and ll<237) then grbp<="010";
	end if;
	if (cc>178 and cc<182 and ll>227 and ll<255) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>245 and ll<255) then grbp<="010";
	end if;
	if (cc>183 and cc<187 and ll>227 and ll<273) then grbp<="010";
	end if;
	if (cc>178 and cc<187 and ll>263 and ll<273) then grbp<="010";
	end if;
end if;

end if;	

-------------------------------mode="111"--------------------tetris---------------------
if mode="111" then

if tstatus/=dead then

	if cc>76 and cc<125 and ll>54 and ll<399 then                
		tccc<=(to_integer(unsigned(cc))-77)/4;
		tlll<=(to_integer(unsigned(ll))-55)/8;                       ------------------39
		if ttstatus1(tccc,tlll)='0' and ttstatus0(tccc,tlll)='1' then
			grbp<="010";
		end if;
		if ttstatus1(tccc,tlll)='1' and ttstatus0(tccc,tlll)='0' then
			grbp<="101";
		end if;
		if ttstatus1(tccc,tlll)='1' and ttstatus0(tccc,tlll)='1' then
			grbp<="111";
		end if;
		if ttstatus1(tccc,tlll)='0' and ttstatus0(tccc,tlll)='0' then
			grbp<="000";
		end if;
	end if;

----------------------------tetris---begin------------------------

	if (cc=162 and ll=78) then grbp<="010";
	end if;
	if (ll=78 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=79 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=80 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=80 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=81 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=81 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=82 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=82 and cc>=149 and cc<151) then grbp<="010";
	end if;
	if (ll=82 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=83 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=83 and cc>=149 and cc<151) then grbp<="010";
	end if;
	if (ll=83 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=84 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=84 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=84 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=85 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (ll=85 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=86 and cc>=129 and cc<137) then grbp<="010";
	end if;
	if (cc=148 and ll=86) then grbp<="010";
	end if;
	if (ll=86 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (cc=169 and ll=86) then grbp<="010";
	end if;
	if (cc=132 and ll=87) then grbp<="010";
	end if;
	if (ll=87 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=87 and cc>=140 and cc<143) then grbp<="010";
	end if;
	if (ll=87 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=87 and cc>=154 and cc<156) then grbp<="010";
	end if;
	if (ll=87 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=87 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=87 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=87) then grbp<="010";
	end if;
	if (cc=132 and ll=88) then grbp<="010";
	end if;
	if (ll=88 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=88 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=88 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=88 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=88 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=88 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=88 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=88) then grbp<="010";
	end if;
	if (ll=88 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=89 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=89 and cc>=139 and cc<144) then grbp<="010";
	end if;
	if (ll=89 and cc>=147 and cc<153) then grbp<="010";
	end if;
	if (ll=89 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=89 and cc>=158 and cc<160) then grbp<="010";
	end if;
	if (ll=89 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=89 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=89) then grbp<="010";
	end if;
	if (ll=89 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=90 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=90 and cc>=138 and cc<145) then grbp<="010";
	end if;
	if (ll=90 and cc>=147 and cc<153) then grbp<="010";
	end if;
	if (ll=90 and cc>=154 and cc<160) then grbp<="010";
	end if;
	if (ll=90 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=90 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=90) then grbp<="010";
	end if;
	if (ll=90 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=91 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=91 and cc>=138 and cc<145) then grbp<="010";
	end if;
	if (ll=91 and cc>=147 and cc<153) then grbp<="010";
	end if;
	if (ll=91 and cc>=154 and cc<160) then grbp<="010";
	end if;
	if (ll=91 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=91 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=91) then grbp<="010";
	end if;
	if (ll=91 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=92 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=92 and cc>=138 and cc<141) then grbp<="010";
	end if;
	if (ll=92 and cc>=142 and cc<145) then grbp<="010";
	end if;
	if (ll=92 and cc>=147 and cc<153) then grbp<="010";
	end if;
	if (ll=92 and cc>=154 and cc<160) then grbp<="010";
	end if;
	if (ll=92 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=92 and cc>=167 and cc<169) then grbp<="010";
	end if;
	if (cc=132 and ll=93) then grbp<="010";
	end if;
	if (ll=93 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=93 and cc>=138 and cc<141) then grbp<="010";
	end if;
	if (ll=93 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (ll=93 and cc>=147 and cc<153) then grbp<="010";
	end if;
	if (ll=93 and cc>=154 and cc<160) then grbp<="010";
	end if;
	if (ll=93 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=93 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=94 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=94 and cc>=138 and cc<140) then grbp<="010";
	end if;
	if (ll=94 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (ll=94 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=94 and cc>=154 and cc<160) then grbp<="010";
	end if;
	if (ll=94 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=94 and cc>=166 and cc<169) then grbp<="010";
	end if;
	if (ll=95 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=95 and cc>=137 and cc<140) then grbp<="010";
	end if;
	if (ll=95 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (ll=95 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=95 and cc>=154 and cc<158) then grbp<="010";
	end if;
	if (ll=95 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=95 and cc>=166 and cc<170) then grbp<="010";
	end if;
	if (ll=96 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=96 and cc>=137 and cc<140) then grbp<="010";
	end if;
	if (ll=96 and cc>=143 and cc<145) then grbp<="010";
	end if;
	if (ll=96 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=96 and cc>=154 and cc<158) then grbp<="010";
	end if;
	if (ll=96 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=96 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=132 and ll=97) then grbp<="010";
	end if;
	if (ll=97 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=97 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=97 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=97 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=97 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=97 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=132 and ll=98) then grbp<="010";
	end if;
	if (ll=98 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=98 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=98 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=98 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=98 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=98 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=98) then grbp<="010";
	end if;
	if (cc=132 and ll=99) then grbp<="010";
	end if;
	if (ll=99 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=99 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=99 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=99 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=99 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=99 and cc>=167 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=99) then grbp<="010";
	end if;
	if (cc=132 and ll=100) then grbp<="010";
	end if;
	if (ll=100 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=100 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=100 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=100 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=100 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=100 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=100) then grbp<="010";
	end if;
	if (ll=100 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=101 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=101 and cc>=137 and cc<145) then grbp<="010";
	end if;
	if (ll=101 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=101 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=101 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=101 and cc>=168 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=101) then grbp<="010";
	end if;
	if (ll=101 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=102 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=102 and cc>=137 and cc<140) then grbp<="010";
	end if;
	if (ll=102 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=102 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=102 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=102 and cc>=169 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=102) then grbp<="010";
	end if;
	if (ll=102 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=103 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=103 and cc>=137 and cc<140) then grbp<="010";
	end if;
	if (ll=103 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=103 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=103 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=103 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=104 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=104 and cc>=137 and cc<140) then grbp<="010";
	end if;
	if (ll=104 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=104 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=104 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=104 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=105 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=105 and cc>=138 and cc<140) then grbp<="010";
	end if;
	if (ll=105 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (ll=105 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=105 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=105 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=106 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=106 and cc>=138 and cc<141) then grbp<="010";
	end if;
	if (cc=148 and ll=106) then grbp<="010";
	end if;
	if (ll=106 and cc>=148 and cc<151) then grbp<="010";
	end if;
	if (cc=154 and ll=106) then grbp<="010";
	end if;
	if (ll=106 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=106 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=106 and cc>=166 and cc<168) then grbp<="010";
	end if;
	if (ll=106 and cc>=170 and cc<173) then grbp<="010";
	end if;
	if (ll=107 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=107 and cc>=138 and cc<145) then grbp<="010";
	end if;
	if (ll=107 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=107 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=107 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=107 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=107) then grbp<="010";
	end if;
	if (ll=107 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=108 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=108 and cc>=138 and cc<145) then grbp<="010";
	end if;
	if (ll=108 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=108 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=108 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=108 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=108) then grbp<="010";
	end if;
	if (ll=108 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=109 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=109 and cc>=138 and cc<145) then grbp<="010";
	end if;
	if (ll=109 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=109 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=109 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=109 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=109) then grbp<="010";
	end if;
	if (ll=109 and cc>=171 and cc<173) then grbp<="010";
	end if;
	if (ll=110 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=110 and cc>=139 and cc<145) then grbp<="010";
	end if;
	if (ll=110 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=110 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=110 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=110 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=110) then grbp<="010";
	end if;
	if (cc=132 and ll=111) then grbp<="010";
	end if;
	if (ll=111 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=111 and cc>=139 and cc<145) then grbp<="010";
	end if;
	if (ll=111 and cc>=148 and cc<153) then grbp<="010";
	end if;
	if (ll=111 and cc>=154 and cc<157) then grbp<="010";
	end if;
	if (ll=111 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=111 and cc>=166 and cc<171) then grbp<="010";
	end if;
	if (cc=171 and ll=111) then grbp<="010";
	end if;
	if (cc=132 and ll=112) then grbp<="010";
	end if;
	if (ll=112 and cc>=132 and cc<135) then grbp<="010";
	end if;
	if (ll=112 and cc>=140 and cc<144) then grbp<="010";
	end if;
	if (ll=112 and cc>=149 and cc<152) then grbp<="010";
	end if;
	if (ll=112 and cc>=155 and cc<157) then grbp<="010";
	end if;
	if (ll=112 and cc>=162 and cc<164) then grbp<="010";
	end if;
	if (ll=112 and cc>=167 and cc<171) then grbp<="010";
	end if;

----------------------------tetris--end------------------------
	
case food0 is                             ------------128-174----135-215-----cc>138+2 and cc<147 and ll>166+4 and ll<183-------------
    when 0=>
    if cc>142 and cc<145 and ll>166 and ll<183 then
		grbp<="011";
	end if;
    when 1=>
    if cc>140 and cc<143 and ll>170 and ll<175 then
		grbp<="011";
	end if;
	if cc>140 and cc<147 and ll>174 and ll<179 then
		grbp<="011";
	end if;
    when 2=>
    if cc>142 and cc<145 and ll>170 and ll<175 then
		grbp<="011";
	end if;
	if cc>140 and cc<147 and ll>174 and ll<179 then
		grbp<="011";
	end if;
    when 3=>
    if cc>144 and cc<147 and ll>170 and ll<175 then
		grbp<="011";
	end if;
	if cc>140 and cc<147 and ll>174 and ll<179 then
		grbp<="011";
	end if;
    when 4=>
    if cc>140 and cc<145 and ll>170 and ll<175 then
		grbp<="011";
	end if;
	if cc>142 and cc<147 and ll>174 and ll<179 then
		grbp<="011";
	end if;
    when 5=>
    if cc>142 and cc<147 and ll>170 and ll<175 then
		grbp<="011";
	end if;
	if cc>140 and cc<145 and ll>174 and ll<179 then
		grbp<="011";
	end if;
    when 6=>
    if cc>140 and cc<145 and ll>170 and ll<179 then
		grbp<="011";
	end if;
end case;

--------------------------score-------begin--------------------

if score1="0001" then
	if (cc>137 and cc<144 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0010" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<138 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0011" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0100" then
	if (cc>130 and cc<138 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0101" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>130 and cc<138 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0110" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>130 and cc<138 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score1="0111" then
	if (cc>130 and cc<138 and ll>225 and ll<232) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score1="1000" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>130 and cc<138 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score1="1001" then
	if (cc>130 and cc<151 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>130 and cc<138 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>143 and cc<151 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>130 and cc<151 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;


if score0="0000" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>152 and cc<159 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>166 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0001" then
	if (cc>159 and cc<166 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0010" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<160 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0011" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0100" then
	if (cc>152 and cc<160 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0101" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>152 and cc<160 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0110" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>152 and cc<160 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>249 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="0111" then
	if (cc>152 and cc<160 and ll>225 and ll<232) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
end if;
if score0="1000" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>152 and cc<160 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;
if score0="1001" then
	if (cc>152 and cc<173 and ll>225 and ll<238) then grbp<="010";
	end if;
	if (cc>152 and cc<160 and ll>225 and ll<262) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>249 and ll<262) then grbp<="010";
	end if;
	if (cc>165 and cc<173 and ll>225 and ll<286) then grbp<="010";
	end if;
	if (cc>152 and cc<173 and ll>273 and ll<286) then grbp<="010";
	end if;
end if;


if PT2="0000" then
	if (cc>128 and cc<139 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>128 and cc<132 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>135 and cc<139 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT2="0001" then
	if (cc>131 and cc<136 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT2="0010" then
	if (cc>128 and cc<139 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>135 and cc<139 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>128 and cc<132 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT2="0011" then
	if (cc>128 and cc<139 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>135 and cc<139 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT2="0100" then
	if (cc>128 and cc<132 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>135 and cc<139 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT2="0101" then
	if (cc>128 and cc<139 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>128 and cc<132 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>135 and cc<139 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>128 and cc<139 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;

if PT3="0000" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0001" then
	if (cc>142 and cc<147 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0010" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0011" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0100" then
	if (cc>139 and cc<143 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0101" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0110" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="0111" then
	if (cc>139 and cc<143 and ll>315 and ll<320) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="1000" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT3="1001" then
	if (cc>139 and cc<150 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>139 and cc<143 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>146 and cc<150 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>139 and cc<150 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;

	IF CC >150 and cc<153 AND ((LL <328 AND LL > 323) or (ll<348 and ll>343)) THEN GRBP <= "111";
	END IF;

if PT4="0000" then
	if (cc>153 and cc<164 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>153 and cc<157 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>160 and cc<164 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT4="0001" then
	if (cc>156 and cc<161 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT4="0010" then
	if (cc>153 and cc<164 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>160 and cc<164 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>153 and cc<157 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT4="0011" then
	if (cc>153 and cc<164 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>160 and cc<164 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT4="0100" then
	if (cc>153 and cc<157 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>160 and cc<164 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT4="0101" then
	if (cc>153 and cc<164 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>153 and cc<157 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>160 and cc<164 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>153 and cc<164 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;

if PT5="0000" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0001" then
	if (cc>167 and cc<172 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0010" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0011" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0100" then
	if (cc>164 and cc<168 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0101" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0110" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>331 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="0111" then
	if (cc>164 and cc<168 and ll>315 and ll<320) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="1000" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;
if PT5="1001" then
	if (cc>164 and cc<175 and ll>315 and ll<324) then grbp<="011";
	end if;
	if (cc>164 and cc<168 and ll>315 and ll<340) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>331 and ll<340) then grbp<="011";
	end if;
	if (cc>171 and cc<175 and ll>315 and ll<356) then grbp<="011";
	end if;
	if (cc>164 and cc<175 and ll>347 and ll<356) then grbp<="011";
	end if;
end if;

end if;

end if;
------------------------------------------mode-logo------------------------------------

if mode="000" then
    
	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=204 and ll=52) then grbp<="001";
	end if;
	if (cc=207 and ll=52) then grbp<="001";
	end if;
	if (cc=219 and ll=52) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=53) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=56 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=57 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=203 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=58 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=203 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=59 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (ll=59 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=59 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=215 and cc<219) then grbp<="001";
	end if;
	if (ll=60 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (cc=204 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (ll=61 and cc>=214 and cc<216) then grbp<="001";
	end if;
	if (cc=220 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=227 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (cc=204 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (ll=62 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=62 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=217 and ll=62) then grbp<="001";
	end if;
	if (cc=220 and ll=62) then grbp<="001";
	end if;
	if (cc=223 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (cc=205 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=63) then grbp<="001";
	end if;
	if (cc=214 and ll=63) then grbp<="001";
	end if;
	if (cc=217 and ll=63) then grbp<="001";
	end if;
	if (cc=220 and ll=63) then grbp<="001";
	end if;
	if (cc=223 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (cc=204 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=212 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=65) then grbp<="001";
	end if;
	if (cc=212 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=66) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=217 and ll=66) then grbp<="001";
	end if;
	if (cc=219 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=202 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=67 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=217 and ll=67) then grbp<="001";
	end if;
	if (cc=219 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=202 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=202 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (ll=69 and cc>=207 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=208 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=70 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=70) then grbp<="001";
	end if;
	if (cc=222 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=208 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=72 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=209 and ll=73) then grbp<="001";
	end if;
	if (cc=220 and ll=73) then grbp<="001";
	end if;
	if (cc=201 and ll=77) then grbp<="001";
	end if;
	if (ll=77 and cc>=201 and cc<229) then grbp<="001";
	end if;
	if (cc=201 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=201 and cc<229) then grbp<="001";
	end if;

	if (cc=204 and ll=51) then grbp<="011";
	end if;
	if (cc=207 and ll=51) then grbp<="011";
	end if;
	if (ll=51 and cc>=207 and cc<209) then grbp<="011";
	end if;
	if (cc=203 and ll=52) then grbp<="011";
	end if;
	if (cc=208 and ll=52) then grbp<="011";
	end if;
	if (cc=219 and ll=53) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=206 and ll=54) then grbp<="011";
	end if;
	if (cc=227 and ll=57) then grbp<="011";
	end if;
	if (cc=216 and ll=58) then grbp<="011";
	end if;
	if (cc=205 and ll=59) then grbp<="011";
	end if;
	if (cc=223 and ll=59) then grbp<="011";
	end if;
	if (cc=207 and ll=60) then grbp<="011";
	end if;
	if (cc=214 and ll=60) then grbp<="011";
	end if;
	if (cc=220 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=203 and ll=61) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=218 and ll=61) then grbp<="011";
	end if;
	if (cc=222 and ll=61) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=203 and ll=62) then grbp<="011";
	end if;
	if (cc=203 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=203 and cc<205) then grbp<="011";
	end if;
	if (cc=219 and ll=63) then grbp<="011";
	end if;
	if (cc=203 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=65) then grbp<="011";
	end if;
	if (cc=214 and ll=65) then grbp<="011";
	end if;
	if (cc=207 and ll=66) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=220 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=220 and cc<224) then grbp<="011";
	end if;
	if (ll=70 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=215 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<204) then grbp<="111";
	end if;
	if (ll=51 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=51 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=51 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=52 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=52 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=52 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=220 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=56 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=57 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=208 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=58) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=59 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=59 and cc>=224 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=224 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=61 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (cc=216 and ll=61) then grbp<="111";
	end if;
	if (cc=219 and ll=61) then grbp<="111";
	end if;
	if (cc=224 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=210 and ll=62) then grbp<="111";
	end if;
	if (cc=213 and ll=62) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (ll=62 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=62 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=62 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=221 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=63 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=64 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=65) then grbp<="111";
	end if;
	if (cc=209 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=220 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=220 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=209 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=209 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=209 and ll=70) then grbp<="111";
	end if;
	if (cc=212 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (ll=71 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=71 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=72 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<209) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (ll=73 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (cc=229 and ll=77) then grbp<="111";
	end if;
	if (cc=200 and ll=78) then grbp<="111";
	end if;
	if (cc=229 and ll=78) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="001" then
    


	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=61 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=226 and ll=52) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=229 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=204 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=223 and ll=71) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (ll=73 and cc>=223 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=65 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=226 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (cc=228 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (cc=228 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="010" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=226 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=228 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=227 and ll=65) then grbp<="011";
	end if;
	if (ll=66 and cc>=227 and cc<229) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=225 and ll=70) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="011" then
    


	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=65) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (ll=66 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=223 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=228 and ll=52) then grbp<="011";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=227 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=226 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=226 and cc<229) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=68 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=59) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=60) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=229 and ll=66) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="100" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=215 and ll=58) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=221 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (cc=213 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=61) then grbp<="001";
	end if;
	if (cc=224 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=224 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=63 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=223 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=223 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=223 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=217 and ll=52) then grbp<="011";
	end if;
	if (cc=204 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=54) then grbp<="011";
	end if;
	if (cc=225 and ll=54) then grbp<="011";
	end if;
	if (ll=54 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=205 and ll=56) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=228 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (cc=218 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=206 and ll=64) then grbp<="011";
	end if;
	if (cc=228 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=210 and ll=67) then grbp<="011";
	end if;
	if (cc=213 and ll=67) then grbp<="011";
	end if;
	if (cc=223 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=69) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=224 and ll=70) then grbp<="011";
	end if;
	if (cc=212 and ll=71) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=226 and ll=72) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=223 and ll=60) then grbp<="111";
	end if;
	if (cc=228 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (cc=226 and ll=61) then grbp<="111";
	end if;
	if (cc=229 and ll=61) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=62 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (ll=67 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=224 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=227 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=227 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;
end if;	

if mode="101" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=226 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=228 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=224 and ll=63) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=224 and ll=66) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=227 and ll=53) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=224 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=225 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=67) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=227 and ll=71) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=56 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=57 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=58 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

if mode="111" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=229 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=211 and ll=68) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=227 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=228 and ll=54) then grbp<="011";
	end if;
	if (cc=217 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=220 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=62 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=224 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=225 and ll=64) then grbp<="011";
	end if;
	if (cc=227 and ll=64) then grbp<="011";
	end if;
	if (cc=206 and ll=65) then grbp<="011";
	end if;
	if (cc=218 and ll=65) then grbp<="011";
	end if;
	if (cc=202 and ll=66) then grbp<="011";
	end if;
	if (cc=210 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=211 and ll=69) then grbp<="011";
	end if;
	if (ll=69 and cc>=211 and cc<213) then grbp<="011";
	end if;
	if (cc=222 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (cc=226 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=228 and ll=78) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=229 and ll=63) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=226 and ll=64) then grbp<="111";
	end if;
	if (cc=229 and ll=64) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=225 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=70 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;

end if;
if mode="110" then
	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (cc=217 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=205 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=227 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=210 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (cc=219 and ll=61) then grbp<="001";
	end if;
	if (cc=221 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=218 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=226 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=210 and ll=67) then grbp<="001";
	end if;
	if (cc=212 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=215 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (cc=218 and ll=70) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=71 and cc>=212 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=73) then grbp<="001";
	end if;
	if (cc=204 and ll=73) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=213 and ll=73) then grbp<="001";
	end if;
	if (cc=215 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=207 and ll=54) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=227 and ll=56) then grbp<="011";
	end if;
	if (cc=209 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=220 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=220 and cc<222) then grbp<="011";
	end if;
	if (cc=213 and ll=60) then grbp<="011";
	end if;
	if (cc=222 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=204 and ll=61) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (cc=214 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=62) then grbp<="011";
	end if;
	if (cc=218 and ll=62) then grbp<="011";
	end if;
	if (cc=221 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="011";
	end if;
	if (cc=221 and ll=63) then grbp<="011";
	end if;
	if (cc=226 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=213 and ll=65) then grbp<="011";
	end if;
	if (cc=222 and ll=65) then grbp<="011";
	end if;
	if (cc=210 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=67) then grbp<="011";
	end if;
	if (cc=224 and ll=68) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=213 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=210 and ll=71) then grbp<="011";
	end if;
	if (cc=221 and ll=71) then grbp<="011";
	end if;
	if (cc=204 and ll=72) then grbp<="011";
	end if;
	if (cc=212 and ll=72) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (cc=207 and ll=73) then grbp<="011";
	end if;
	if (cc=209 and ll=73) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;
	if (cc=218 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=223 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=51 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=54 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (cc=217 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=217 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (cc=223 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=63 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=64 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=65 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=66 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=222 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=216 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=205 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

end process;

hs<=hs1;vs<=vs1;r<=grb(2);g<=grb(3);b<=grb(1);

end one;
