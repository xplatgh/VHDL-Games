library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity bigbang is
port(
	clk,rst : in std_logic;
	rxd : in std_logic;
	hs,vs,r,g,b : out std_logic);
end bigbang;

architecture one of bigbang is

signal hs1,vs1,fclk,cclk,sclk,md : std_logic;
signal fs : std_logic_vector(2 downto 0);
signal cc : std_logic_vector(8 downto 0);
signal ll : std_logic_vector(8 downto 0);
signal grbx : std_logic_vector(3 downto 1);
signal grby : std_logic_vector(3 downto 1);
signal grbp : std_logic_vector(3 downto 1);
signal grb : std_logic_vector(3 downto 1);
signal grbc : std_logic_vector(3 downto 1);
signal mode : std_logic_vector(2 downto 0);

signal clk_cnt,clk_rsclk : std_logic_vector(24 downto 0);
signal PT0,PT1,PT2,PT3,PT4,PT5 : std_logic_vector(3 downto 0);
signal pt : std_logic;

signal freq,scal, sin,tri,squ,rl : std_logic;
type index_type is array(0 to 800) of integer range 0 to 200;
signal tri_ind,squ_ind,sin_ind,sin_id : index_type;
signal x : integer range 0 to 200;
signal sin_y,tri_y,squ_y : integer range 0 to 200;
signal wi : integer range 0 to 7;
signal f,sc : integer range 1 to 8;
signal cci : integer range 0 to 511;
signal rrll : integer range 0 to 200;
signal xt : integer range 0 to 1800;

signal clk_rscnt:integer range 0 to 651;
signal sam_clk:std_logic;
type status_type is(start,data,over);
signal status:status_type;
signal sam_cnt:std_logic_vector(2 downto 0);
signal bit_cnt:std_logic_vector(3 downto 0);
signal rcv_shift_reg:std_logic_vector(7 downto 0);
signal rcv_data:std_logiC_vector(7 downto 0);
signal rrr,l,rot,rev,speed,pul : std_logic;
signal rrrr,uu,lll,dd : std_logic;

type status_stype is array(0 to 11,0 to 11) of std_logic;    --(250-2*2)*(400-4*2)/8=12054--------------64x64--------------
type index_stype is array(0 to 100) of integer range 0 to 127;       --max : 12054--------------4096-------
signal status1,status0 : status_stype;
signal index_x,index_y : index_stype;
signal alive : std_logic;
signal di,dir : std_logic_vector(1 downto 0);
signal k : integer range 0 to 127;
signal len : integer range 0 to 100;
signal food : std_logic;
signal food_x,food_y,fx_cnt,fy_cnt : integer range 1 to 10;
signal lcx : std_logic;
signal score1,score0 : std_logic_vector(3 downto 0);
signal ccc,llc : integer range 0 to 127;

type ttstatus_type is array(0 to 11,0 to 42) of std_logic;    --(250-2*2)*(400-4*2)/8=12054
type index_typex is array(0 to 3) of integer range 0 to 15;
type index_typey is array(0 to 3) of integer range 0 to 63;
type tstatuse_type is (start,usual,dead);
signal ttstatus1,ttstatus0 : ttstatus_type;
signal tindex_x : index_typex;
signal tindex_y : index_typey;
signal tstatus : tstatuse_type;
signal food0,food1,food_cnt : integer range 0 to 6;
signal tra,tra_r,tra_l,tra_ro,tra_re,tra_d : std_logic;
signal ti,tj,tk,tm,tn,tsp : integer range 0 to 63;
signal tccc,tlll : integer range 0 to 511;

begin
grb(2)<=(grbp(2))and hs1 and vs1;
grb(3)<=(grbp(3))and hs1 and vs1;
grb(1)<=(grbp(1))and hs1 and vs1;


------------------------------------rs232-------------------------------

P1:process(clk,rst)
begin
	if rst='0' then
		clk_rscnt<=0;
	elsif rising_edge(clk) then
		if clk_rscnt=651 then
			clk_rscnt<=0;
			sam_clk<='1';
		else
			clk_rscnt<=clk_rscnt+1;
			sam_clk<='0';
		end if;
	end if;
end process P1;

P2:process(clk,rst)
begin
	if rst='0' then
		status<=start;
		sam_cnt<="000";
		bit_cnt<="0000";
		rcv_shift_reg<="00111111";
		rcv_data<="00111111";

		freq<='0';
		scal<='0'; 
		sin<='1';
		tri<='1';
		squ<='1';
		rl<='0';
		rrll<=0;

		rrr<='0';
		l<='0';
		rot<='0';
		rev<='0';
		speed<='0';
		pul<='0';

		rrrr<='0';
		uu<='0';
		lll<='0';
		dd<='0';

	elsif rising_edge(clk) then
		if sam_clk='1' then
			case status is
				when start=>
					if rxd='0' then
						if sam_cnt="011" then
							sam_cnt<="000";
							status<=data;
							bit_cnt<="0000";
						else
							sam_cnt<=sam_cnt+'1';
						end if;
					end if;
				when data=>
					if sam_cnt="111" then
						if bit_cnt="1000" then
							status<=over;
						else
							rcv_shift_reg<=rxd&rcv_shift_reg(7 downto 1);
							sam_cnt<="000";
							bit_cnt<=bit_cnt+'1';
						end if;
					else
						sam_cnt<=sam_cnt+'1';
					end if;
				when over=>
					rcv_data<=rcv_shift_reg;
					
					if rcv_data="00001010" then
						if mode="111" then               
							mode<="000";
						else
							mode<=mode+1;
						end if;		
					end if;	
					mode<="110";	
					if mode="101" then
						if rcv_data="01110001" then
							if f=8 then
							f<=1;
							else
							f<=f+1;
							end if;
						elsif rcv_data="01110111" then
							if sc=8 then
							sc<=1;
							elsif (sc=1 or sc=2 or sc=4) then
							sc<=sc*2;
							else
							sc<=1;
							end if;
						elsif rcv_data="01100101" then
							sin<=not sin;
						elsif rcv_data="01110010" then
							tri<=not tri;
						elsif rcv_data="01110100" then
							squ<=not squ;
						elsif rcv_data="01111001" then
							if rrll=200 then
							rrll<=0;
							else 
							rrll<=rrll+1;
							end if;
						end if;	
								
					elsif mode="111" then
						if rcv_data="01100001" then
							rrr<=not rrr;
						elsif rcv_data="01110011" then
							l<=not l;
						elsif rcv_data="01100100" then
							rot<=not rot;
						elsif rcv_data="01100110" then
							rev<=not rev;
						elsif rcv_data="01100111" then
							speed<=not speed;
						elsif rcv_data="01101000" then
							pul<=not pul;
						end if;
					elsif mode="110" then
						if rcv_data="01111010" then
							rrrr<=not rrrr;
						elsif rcv_data="01111000" then
							uu<=not uu;
						elsif rcv_data="01100011" then
							lll<=not lll;
						elsif rcv_data="01110110" then
							dd<=not dd;
						end if;
					end if;
					
					status<=start;
			end case;
		end if;
	end if;
end process P2;


    PROCESS( CLK )
    BEGIN
        IF CLK'EVENT AND CLK = '1' THEN -- 50MHz 5分频
            IF FS = 4 THEN FS <= "000";
            ELSE
                FS <= (FS + 1);
            END IF;
        END IF;
    END PROCESS;
    FCLK <= FS(2);
    PROCESS( FCLK )--再315分频，12000000/(13*30)=30769,接近于行频31469
    BEGIN
        IF FCLK'EVENT AND FCLK = '1' THEN
            IF CC = 314 THEN  CC <= "000000000";
            ELSE
                CC <= CC + 1;
            END IF;
        END IF;
    END PROCESS;
    CCLK <= CC(8);
    
    PROCESS( CCLK )
    BEGIN
        IF CCLK'EVENT AND CCLK = '0' THEN
            IF LL = 481 THEN  LL <= "000000000";
            ELSE
                LL <= LL + 1;
            END IF;
        END IF;
    END PROCESS;
    
    
    PROCESS( CC,LL )
    BEGIN
        IF CC > 251 THEN  HS1 <= '0';  --行同步
        ELSE
            HS1 <= '1';
        END IF;
        IF LL > 479 THEN  VS1 <= '0'; --场同步
        ELSE
            VS1 <= '1';
        END IF;
    END PROCESS;
    
process(clk)
begin
	if rising_edge(clk) then
		IF clk_cnt=25000000 THEN clk_cnt<=(others=>'0');
        ELSE
            clk_cnt<=clk_cnt+1;
        END IF;
    END IF;
END PROCESS;

sclk<=clk_cnt(24);
----------------------------------------clk------------------------------
process(sclk,rst)
begin
if rst='0' then

PT0<="0000";PT1<="0000";PT2<="0000";PT3<="0000";PT4<="0000";PT5<="0000";pt<='0';

elsif rising_edge(sclk) then
pt<=not pt;
if pt='1' then
	if PT4="0101" and PT5="1001" then
		if PT2="0101" and PT3="1001" then
			if PT0="0010" and PT1="0011" then
				PT0<="0000";PT1<="0000";
			elsif PT1="1001" then
				PT0<=PT0+1;PT1<="0000";
			else
				PT1<=PT1+1;
			end if;
			PT2<="0000";PT3<="0000";
		elsif PT3="1001" then
			PT2<=PT2+1;PT3<="0000";
		else
			PT3<=PT3+1;
		end if;
		PT4<="0000";PT5<="0000";
	elsif PT5="1001" then
		PT4<=PT4+1;PT5<="0000";
	else
		PT5<=PT5+1;
	end if;
end if;
end if;
end process;

 ------------------------------------------wave---------------------------------   

---------------------snake------------------------

process(clk, rst)
begin

if (rst='0') then
if mode="110" then
	di<="00";    --right 
	for i in 0 to 11 loop 
		for j in 0 to 11 loop
			if (i=0 or i=11 or j=0 or j=11) then
				status1(i,j)<='1';
				status0(i,j)<='1';
			else
				status1(i,j)<='0';           --"00":free;  "01":snake&wall;   "10":food
				status0(i,j)<='0';
			end if;
		end loop;
	end loop;
	status1(6,6)<='0';
	status0(6,6)<='1';
	status1(5,6)<='0';
	status0(5,6)<='1';
	status1(4,6)<='0';
	status0(4,6)<='1';
	index_x(0)<=6;
	index_y(0)<=6;
	index_x(1)<=5;
	index_y(1)<=6;
	index_x(2)<=4;
	index_y(2)<=6;
	for i in 3 to 100 loop
		index_x(i)<=0;
		index_y(i)<=0;
	end loop;
	alive<='1';
	len<=2;
	food<='0';
	food_x<=fx_cnt;
	food_y<=fy_cnt;
	if (status1(food_x,food_y)='0' and status0(food_x,food_y)='0') then
		status1(food_x,food_y)<='1';
		status0(food_x,food_y)<='0';
		food<='1';
	end if; 
end if;
score1<="0000";
score0<="0000";

elsif rising_edge(clk) then

if mode="110" then
if fx_cnt=10 then
	fx_cnt<=1;
else
	fx_cnt<=fx_cnt+1;
end if;
if fy_cnt=1 then
	fy_cnt<=10;
else
	fy_cnt<=fy_cnt-1;
end if;
if fx_cnt+food_x>10 then
	fx_cnt<=fx_cnt+food_x-10;
else
	fx_cnt<=fx_cnt+food_x;
end if;
if fy_cnt>food_y then
	fy_cnt<=fy_cnt-food_y;
else
	fy_cnt<=fy_cnt+10-food_y;
end if;

if rrrr='1' then
	dir<="00";
elsif uu='1' then
	dir<="01";
elsif lll='1' then
	dir<="10";
elsif dd='1' then
	dir<="11";
else
	dir<="00";
end if;
end if;

if lcx='0' and sclk='1' then

if mode="110" then

if fx_cnt=10 then
	fx_cnt<=1;
else
	fx_cnt<=fx_cnt+1;
end if;
if fy_cnt=1 then
	fy_cnt<=10;
else
	fy_cnt<=fy_cnt-1;
end if;

	if (di(0) xor dir(0))='1' then
		di<=dir;
	end if;	
	status1(index_x(0),index_y(0))<='0';
	status0(index_x(0),index_y(0))<='1';
	status1(index_x(len+1),index_y(len+1))<='0';
	status0(index_x(len+1),index_y(len+1))<='0';
	if (di="00" and alive='1') then        --right
		if  status0(index_x(0)+1,index_y(0))='1' then
			alive<='0';
		elsif status1(index_x(0)+1,index_y(0))='1' and status0(index_x(0)+1,index_y(0))='0' then
			food<='0';
			if (len<99) then
				len<=len+1;
			end if;
			if score1="1001" and score0="1001" then
				score1<="0000";
				score0<="0000";
			elsif score0="1001" then
				score1<=score1+1;
				score0<="0000";
			else
				score0<=score0+1;
			end if;
		end if;
		for k in 0 to 99 loop
			if k<=len then
				index_x(k+1)<=index_x(k);
				index_y(k+1)<=index_y(k);
			end if;
		end loop;
		index_x(0)<=index_x(0)+1;
	elsif (di="01" and alive='1') then    --up
		if  status0(index_x(0),index_y(0)-1)='1' then
			alive<='0';
		elsif status1(index_x(0),index_y(0)-1)='1' and status0(index_x(0),index_y(0)-1)='0' then
			food<='0';
			if (len<99) then
				len<=len+1;
			end if;
			if score1="1001" and score0="1001" then
				score1<="0000";
				score0<="0000";
			elsif score0="1001" then
				score1<=score1+1;
				score0<="0000";
			else
				score0<=score0+1;
			end if;
		else
		for k in 0 to 99 loop
			if k<=len then
				index_x(k+1)<=index_x(k);
				index_y(k+1)<=index_y(k);
			end if;
		end loop;
		index_y(0)<=index_y(0)-1;
		end if;
	elsif (di="10" and alive='1') then    --left
		if status0(index_x(0)-1,index_y(0))='1' then
			alive<='0';
		elsif status1(index_x(0)-1,index_y(0))='1' and status0(index_x(0)-1,index_y(0))='0' then
			food<='0';
			if (len<99) then
				len<=len+1;
			end if;
			if score1="1001" and score0="1001" then
				score1<="0000";
				score0<="0000";
			elsif score0="1001" then
				score1<=score1+1;
				score0<="0000";
			else
				score0<=score0+1;
			end if;
		else
		for k in 0 to 99 loop
			if k<=len then
				index_x(k+1)<=index_x(k);
				index_y(k+1)<=index_y(k);
			end if;
		end loop;
		index_x(0)<=index_x(0)-1;
		end if;
	elsif (di="11" and alive='1') then    --down
		if  status0(index_x(0),index_y(0)+1)='1' then
			alive<='0';
		elsif status1(index_x(0),index_y(0)+1)='1' and status0(index_x(0),index_y(0)+1)='0' then
			food<='0';
			if (len<99) then
				len<=len+1;
			end if;
			if score1="1001" and score0="1001" then
				score1<="0000";
				score0<="0000";
			elsif score0="1001" then
				score1<=score1+1;
				score0<="0000";
			else
				score0<=score0+1;
			end if;
		else
		for k in 0 to 99 loop
			if k<=len then
				index_x(k+1)<=index_x(k);
				index_y(k+1)<=index_y(k);
			end if;
		end loop;
		index_y(0)<=index_y(0)+1;	
		end if;
	end if;

if alive='1' and food='0' then
	food_x<=fx_cnt;
	food_y<=fy_cnt;
	if (status1(food_x,food_y)='0' and status0(food_x,food_y)='0') then
		status1(food_x,food_y)<='1';
		status0(food_x,food_y)<='0';
		food<='1';
	end if;
end if;
status1(0,0)<='1';status0(0,0)<='1';
end if;	
-------------------------------tetris------------------------

end if;	
lcx<=sclk;
end if;	

end process;
				
process(cc,ll)
begin 
	grbp<="000";


--------------------------------mode="000"--------------------vertical--------------------

-------------------------------mode="110"--------------------snake---------------------
if mode="110" and alive='1' then
	 if cc>89 and cc<137 and ll>100 and ll<195 then
	 ccc<=to_integer(unsigned(cc-90))/4;
	 llc<=to_integer(unsigned(ll-100))/8;

	if status1(ccc,llc)='1' and status0(ccc,llc)='1' then
		grbp<="010";
	elsif status1(ccc,llc)='0' and status0(ccc,llc)='1' then
		grbp<="101";
	elsif status1(ccc,llc)='1' and status0(ccc,llc)='0' then
		grbp<="011";
	end if;
	 end if;
	----------------------------------snake---------begin----------------------

	if (cc=60 and ll=337) then grbp<="010";
	end if;
	if (ll=337 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=338 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=339 and cc>=38 and cc<40) then grbp<="010";
	end if;
	if (ll=339 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=340 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (ll=340 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=341 and cc>=37 and cc<42) then grbp<="010";
	end if;
	if (ll=341 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=342 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=342 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=343 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=343 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=344 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=344 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=345 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=345 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=346 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (cc=54 and ll=346) then grbp<="010";
	end if;
	if (ll=346 and cc>=54 and cc<56) then grbp<="010";
	end if;
	if (ll=346 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=346 and cc>=70 and cc<72) then grbp<="010";
	end if;
	if (cc=36 and ll=347) then grbp<="010";
	end if;
	if (ll=347 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=347 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=347 and cc>=46 and cc<49) then grbp<="010";
	end if;
	if (ll=347 and cc>=53 and cc<57) then grbp<="010";
	end if;
	if (ll=347 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=347 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=347 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=347) then grbp<="010";
	end if;
	if (cc=36 and ll=348) then grbp<="010";
	end if;
	if (ll=348 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=348 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=348 and cc>=46 and cc<49) then grbp<="010";
	end if;
	if (ll=348 and cc>=52 and cc<57) then grbp<="010";
	end if;
	if (ll=348 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=348 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=348 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=348) then grbp<="010";
	end if;
	if (cc=36 and ll=349) then grbp<="010";
	end if;
	if (ll=349 and cc>=36 and cc<38) then grbp<="010";
	end if;
	if (ll=349 and cc>=43 and cc<45) then grbp<="010";
	end if;
	if (ll=349 and cc>=46 and cc<50) then grbp<="010";
	end if;
	if (ll=349 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=349 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=349 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=349 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=349) then grbp<="010";
	end if;
	if (cc=36 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=36 and cc<39) then grbp<="010";
	end if;
	if (ll=350 and cc>=43 and cc<50) then grbp<="010";
	end if;
	if (ll=350 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=350 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=350 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=350 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=350) then grbp<="010";
	end if;
	if (ll=350 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=351 and cc>=36 and cc<39) then grbp<="010";
	end if;
	if (ll=351 and cc>=43 and cc<50) then grbp<="010";
	end if;
	if (ll=351 and cc>=53 and cc<58) then grbp<="010";
	end if;
	if (ll=351 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=351 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=351 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=351) then grbp<="010";
	end if;
	if (ll=351 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=352 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=352 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=352 and cc>=47 and cc<50) then grbp<="010";
	end if;
	if (cc=55 and ll=352) then grbp<="010";
	end if;
	if (ll=352 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=352 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=352 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=352 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=352 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=353 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=353 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=353 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=353 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=353 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=353 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (ll=353 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=353 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=354 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=354 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=354 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=354 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=354 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=354 and cc>=63 and cc<65) then grbp<="010";
	end if;
	if (ll=354 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=354 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=355 and cc>=37 and cc<41) then grbp<="010";
	end if;
	if (ll=355 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=355 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=355 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=355 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=355 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=355 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=356 and cc>=37 and cc<42) then grbp<="010";
	end if;
	if (ll=356 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=356 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=356 and cc>=53 and cc<58) then grbp<="010";
	end if;
	if (ll=356 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=356 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=356) then grbp<="010";
	end if;
	if (ll=356 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=357 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (ll=357 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=357 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=357 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=357 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=357 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=357) then grbp<="010";
	end if;
	if (ll=357 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=358 and cc>=38 and cc<42) then grbp<="010";
	end if;
	if (ll=358 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=358 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=358 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=358 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=358 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=358) then grbp<="010";
	end if;
	if (ll=358 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=359 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=359 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=359 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=359 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=359 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=359 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=359) then grbp<="010";
	end if;
	if (ll=359 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=360 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=360 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=360 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=360 and cc>=52 and cc<54) then grbp<="010";
	end if;
	if (ll=360 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=360 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=360 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=360) then grbp<="010";
	end if;
	if (ll=360 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=361 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=361 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=361 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=361 and cc>=52 and cc<54) then grbp<="010";
	end if;
	if (ll=361 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=361 and cc>=60 and cc<65) then grbp<="010";
	end if;
	if (ll=361 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=362 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=362 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=362 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=362 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=362 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=362 and cc>=60 and cc<66) then grbp<="010";
	end if;
	if (ll=362 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=363 and cc>=40 and cc<42) then grbp<="010";
	end if;
	if (ll=363 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=363 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=363 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=363 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=363 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=363 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=363 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (cc=39 and ll=364) then grbp<="010";
	end if;
	if (ll=364 and cc>=39 and cc<42) then grbp<="010";
	end if;
	if (ll=364 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=364 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=364 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=364 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=364 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=364 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=364 and cc>=68 and cc<70) then grbp<="010";
	end if;
	if (ll=365 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=365 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=365 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=365 and cc>=51 and cc<54) then grbp<="010";
	end if;
	if (ll=365 and cc>=55 and cc<58) then grbp<="010";
	end if;
	if (ll=365 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=365 and cc>=63 and cc<66) then grbp<="010";
	end if;
	if (ll=365 and cc>=68 and cc<71) then grbp<="010";
	end if;
	if (cc=36 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=36 and cc<42) then grbp<="010";
	end if;
	if (ll=366 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=366 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=366 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=366 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=366 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=366 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=366) then grbp<="010";
	end if;
	if (ll=366 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=367 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=367 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=367 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=367 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=367 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=367 and cc>=64 and cc<66) then grbp<="010";
	end if;
	if (ll=367 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=367) then grbp<="010";
	end if;
	if (ll=367 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=368 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=368 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=368 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=368 and cc>=52 and cc<58) then grbp<="010";
	end if;
	if (ll=368 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=368 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=368 and cc>=68 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=368) then grbp<="010";
	end if;
	if (ll=368 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=369 and cc>=36 and cc<41) then grbp<="010";
	end if;
	if (ll=369 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=369 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=369 and cc>=52 and cc<55) then grbp<="010";
	end if;
	if (ll=369 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=369 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=369 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=369 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=369) then grbp<="010";
	end if;
	if (ll=369 and cc>=72 and cc<74) then grbp<="010";
	end if;
	if (ll=370 and cc>=36 and cc<40) then grbp<="010";
	end if;
	if (ll=370 and cc>=43 and cc<46) then grbp<="010";
	end if;
	if (ll=370 and cc>=48 and cc<50) then grbp<="010";
	end if;
	if (ll=370 and cc>=52 and cc<55) then grbp<="010";
	end if;
	if (ll=370 and cc>=56 and cc<58) then grbp<="010";
	end if;
	if (ll=370 and cc>=60 and cc<62) then grbp<="010";
	end if;
	if (ll=370 and cc>=64 and cc<67) then grbp<="010";
	end if;
	if (ll=370 and cc>=69 and cc<72) then grbp<="010";
	end if;
	if (cc=72 and ll=370) then grbp<="010";
	end if;
	if (cc=38 and ll=371) then grbp<="010";
	end if;
	if (cc=53 and ll=371) then grbp<="010";
	end if;
	if (cc=70 and ll=371) then grbp<="010";
	end if;
	if (ll=371 and cc>=70 and cc<72) then grbp<="010";
	end if;


-------------------------------------snake--------------end-------------------

---------------------------------------time-----------begin-------------------

if cc>123 and cc<127 and ll>341 and ll<348 then
	grbp<="010";
end if;
if cc>123 and cc<127 and ll>362 and ll<369 then
	grbp<="010";
end if;

if PT2="0000" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0001" then
	if (cc>95 and cc<101 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0010" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0011" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0100" then
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0101" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0110" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="0111" then
	if (cc>90 and cc<96 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="1000" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT2="1001" then
	if (cc>90 and cc<106 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>90 and cc<96 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>100 and cc<106 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>90 and cc<106 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT3="0000" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0001" then
	if (cc>111 and cc<117 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0010" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0011" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0100" then
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0101" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0110" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="0111" then
	if (cc>106 and cc<112 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="1000" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT3="1001" then
	if (cc>106 and cc<122 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>106 and cc<112 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>116 and cc<122 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>106 and cc<122 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT4="0000" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0001" then
	if (cc>133 and cc<139 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0010" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0011" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0100" then
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0101" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0110" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="0111" then
	if (cc>128 and cc<134 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="1000" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT4="1001" then
	if (cc>128 and cc<144 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>128 and cc<134 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>138 and cc<144 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>128 and cc<144 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if PT5="0000" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0001" then
	if (cc>149 and cc<155 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0010" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0011" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0100" then
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0101" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0110" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="0111" then
	if (cc>144 and cc<150 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="1000" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if PT5="1001" then
	if (cc>144 and cc<160 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>144 and cc<150 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>154 and cc<160 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>144 and cc<160 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;



---------------------------------------time-------------end---------------------

--------------------------------------score--------------begin-----------------

if score1="0000" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<188 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>194 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0001" then
	if (cc>188 and cc<194 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0010" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0011" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0100" then
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0101" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0110" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="0111" then
	if (cc>183 and cc<189 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score1="1000" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score1="1001" then
	if (cc>183 and cc<199 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>183 and cc<189 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>193 and cc<199 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>183 and cc<199 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

if score0="0000" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<204 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>210 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0001" then
	if (cc>204 and cc<210 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0010" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0011" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0100" then
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0101" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0110" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>351 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="0111" then
	if (cc>199 and cc<205 and ll>335 and ll<340) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
end if;
if score0="1000" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;
if score0="1001" then
	if (cc>199 and cc<215 and ll>335 and ll<344) then grbp<="010";
	end if;
	if (cc>199 and cc<205 and ll>335 and ll<360) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>351 and ll<360) then grbp<="010";
	end if;
	if (cc>209 and cc<215 and ll>335 and ll<376) then grbp<="010";
	end if;
	if (cc>199 and cc<215 and ll>367 and ll<376) then grbp<="010";
	end if;
end if;

--------------------------------------score---------end---------------------------


	---------------------------------------------------------------35-75-90-106-122-128-144-160-183-199-215---------
	---------------------------------------------------------------54-318-335-375--------------------------

end if;


------------------------------------------mode-logo------------------------------------

if mode="000" then
    
	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=204 and ll=52) then grbp<="001";
	end if;
	if (cc=207 and ll=52) then grbp<="001";
	end if;
	if (cc=219 and ll=52) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=53) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=56 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=57 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=203 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=58 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=203 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=59 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (ll=59 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=59 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=215 and cc<219) then grbp<="001";
	end if;
	if (ll=60 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (cc=204 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (ll=61 and cc>=214 and cc<216) then grbp<="001";
	end if;
	if (cc=220 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=227 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (cc=204 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (ll=62 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=62 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=217 and ll=62) then grbp<="001";
	end if;
	if (cc=220 and ll=62) then grbp<="001";
	end if;
	if (cc=223 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (cc=205 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=63) then grbp<="001";
	end if;
	if (cc=214 and ll=63) then grbp<="001";
	end if;
	if (cc=217 and ll=63) then grbp<="001";
	end if;
	if (cc=220 and ll=63) then grbp<="001";
	end if;
	if (cc=223 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (cc=204 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=204 and cc<207) then grbp<="001";
	end if;
	if (cc=212 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=212 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=65) then grbp<="001";
	end if;
	if (cc=212 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<224) then grbp<="001";
	end if;
	if (cc=202 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=66) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=217 and ll=66) then grbp<="001";
	end if;
	if (cc=219 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=202 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=67 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=217 and ll=67) then grbp<="001";
	end if;
	if (cc=219 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=202 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=202 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (ll=69 and cc>=207 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=208 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (ll=70 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (cc=219 and ll=70) then grbp<="001";
	end if;
	if (cc=222 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=208 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<211) then grbp<="001";
	end if;
	if (ll=72 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=209 and ll=73) then grbp<="001";
	end if;
	if (cc=220 and ll=73) then grbp<="001";
	end if;
	if (cc=201 and ll=77) then grbp<="001";
	end if;
	if (ll=77 and cc>=201 and cc<229) then grbp<="001";
	end if;
	if (cc=201 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=201 and cc<229) then grbp<="001";
	end if;

	if (cc=204 and ll=51) then grbp<="011";
	end if;
	if (cc=207 and ll=51) then grbp<="011";
	end if;
	if (ll=51 and cc>=207 and cc<209) then grbp<="011";
	end if;
	if (cc=203 and ll=52) then grbp<="011";
	end if;
	if (cc=208 and ll=52) then grbp<="011";
	end if;
	if (cc=219 and ll=53) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=206 and ll=54) then grbp<="011";
	end if;
	if (cc=227 and ll=57) then grbp<="011";
	end if;
	if (cc=216 and ll=58) then grbp<="011";
	end if;
	if (cc=205 and ll=59) then grbp<="011";
	end if;
	if (cc=223 and ll=59) then grbp<="011";
	end if;
	if (cc=207 and ll=60) then grbp<="011";
	end if;
	if (cc=214 and ll=60) then grbp<="011";
	end if;
	if (cc=220 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=203 and ll=61) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=218 and ll=61) then grbp<="011";
	end if;
	if (cc=222 and ll=61) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=203 and ll=62) then grbp<="011";
	end if;
	if (cc=203 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=203 and cc<205) then grbp<="011";
	end if;
	if (cc=219 and ll=63) then grbp<="011";
	end if;
	if (cc=203 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=64) then grbp<="011";
	end if;
	if (cc=211 and ll=65) then grbp<="011";
	end if;
	if (cc=214 and ll=65) then grbp<="011";
	end if;
	if (cc=207 and ll=66) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=220 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=220 and cc<224) then grbp<="011";
	end if;
	if (ll=70 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=215 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<204) then grbp<="111";
	end if;
	if (ll=51 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=51 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=51 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=52 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=52 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=52 and cc>=220 and cc<229) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=220 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=56 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=57 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=208 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=58) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=59 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=59 and cc>=224 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=224 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=61 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (cc=216 and ll=61) then grbp<="111";
	end if;
	if (cc=219 and ll=61) then grbp<="111";
	end if;
	if (cc=224 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=210 and ll=62) then grbp<="111";
	end if;
	if (cc=213 and ll=62) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (ll=62 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=62 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=62 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=221 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=63 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=64 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=65) then grbp<="111";
	end if;
	if (cc=209 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=215 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=224 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<217) then grbp<="111";
	end if;
	if (cc=220 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=220 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=209 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=209 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=209 and ll=70) then grbp<="111";
	end if;
	if (cc=212 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (ll=71 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=71 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=72 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<209) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<214) then grbp<="111";
	end if;
	if (ll=73 and cc>=215 and cc<220) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (cc=229 and ll=77) then grbp<="111";
	end if;
	if (cc=200 and ll=78) then grbp<="111";
	end if;
	if (cc=229 and ll=78) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="001" then
    


	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=61 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=226 and ll=52) then grbp<="011";
	end if;
	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=229 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=66 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=204 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=223 and ll=71) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (ll=73 and cc>=223 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=65 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (ll=68 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=226 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (cc=228 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (cc=228 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="010" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=226 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=64 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=55) then grbp<="011";
	end if;
	if (cc=228 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=228 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=227 and ll=65) then grbp<="011";
	end if;
	if (ll=66 and cc>=227 and cc<229) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=225 and ll=70) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="011" then
    


	if (cc=229 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=229 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=227 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=62 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=65) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (ll=66 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=223 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=223 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=222 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=228 and ll=52) then grbp<="011";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="011";
	end if;
	if (cc=218 and ll=55) then grbp<="011";
	end if;
	if (cc=227 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=215 and ll=58) then grbp<="011";
	end if;
	if (cc=226 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=226 and cc<229) then grbp<="011";
	end if;
	if (ll=64 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=201 and ll=66) then grbp<="011";
	end if;
	if (ll=68 and cc>=201 and cc<203) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=215 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<229) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=59) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (cc=229 and ll=60) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=228 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=64 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=64 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=229 and ll=66) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<226) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;
end if;
if mode="100" then
    


	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=215 and ll=58) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=221 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=211 and ll=61) then grbp<="001";
	end if;
	if (cc=213 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=61) then grbp<="001";
	end if;
	if (cc=224 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=224 and ll=62) then grbp<="001";
	end if;
	if (cc=227 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=63 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=227 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=227 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=227 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=221 and cc<224) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=223 and ll=69) then grbp<="001";
	end if;
	if (cc=226 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=212 and cc<214) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=223 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=223 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=224 and cc<226) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=217 and ll=52) then grbp<="011";
	end if;
	if (cc=204 and ll=53) then grbp<="011";
	end if;
	if (cc=204 and ll=54) then grbp<="011";
	end if;
	if (cc=225 and ll=54) then grbp<="011";
	end if;
	if (ll=54 and cc>=225 and cc<227) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=205 and ll=56) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (ll=61 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=228 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=228 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (cc=218 and ll=63) then grbp<="011";
	end if;
	if (cc=228 and ll=63) then grbp<="011";
	end if;
	if (cc=206 and ll=64) then grbp<="011";
	end if;
	if (cc=228 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=210 and ll=67) then grbp<="011";
	end if;
	if (cc=213 and ll=67) then grbp<="011";
	end if;
	if (cc=223 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=68) then grbp<="011";
	end if;
	if (cc=213 and ll=69) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=219 and ll=70) then grbp<="011";
	end if;
	if (cc=224 and ll=70) then grbp<="011";
	end if;
	if (cc=212 and ll=71) then grbp<="011";
	end if;
	if (cc=218 and ll=72) then grbp<="011";
	end if;
	if (cc=226 and ll=72) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=223 and ll=60) then grbp<="111";
	end if;
	if (cc=228 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (cc=226 and ll=61) then grbp<="111";
	end if;
	if (cc=229 and ll=61) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (ll=62 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<227) then grbp<="111";
	end if;
	if (ll=65 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=66 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<223) then grbp<="111";
	end if;
	if (ll=67 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=67 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=224 and cc<227) then grbp<="111";
	end if;
	if (ll=68 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=224 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=224 and cc<226) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=227 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=227 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=214 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;
end if;	

if mode="101" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (cc=203 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=227 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=226 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=226 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=226 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=59 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=61) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (cc=228 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=219 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=224 and ll=63) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=219 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (cc=224 and ll=66) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=226 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=208 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=227 and ll=53) then grbp<="011";
	end if;
	if (cc=217 and ll=54) then grbp<="011";
	end if;
	if (cc=204 and ll=55) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=210 and ll=58) then grbp<="011";
	end if;
	if (cc=221 and ll=58) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=213 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=214 and ll=62) then grbp<="011";
	end if;
	if (cc=224 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=63) then grbp<="011";
	end if;
	if (cc=217 and ll=63) then grbp<="011";
	end if;
	if (cc=225 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=208 and ll=64) then grbp<="011";
	end if;
	if (cc=218 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=212 and ll=67) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=69) then grbp<="011";
	end if;
	if (cc=222 and ll=69) then grbp<="011";
	end if;
	if (cc=212 and ll=70) then grbp<="011";
	end if;
	if (cc=214 and ll=70) then grbp<="011";
	end if;
	if (cc=227 and ll=71) then grbp<="011";
	end if;
	if (cc=207 and ll=72) then grbp<="011";
	end if;
	if (cc=216 and ll=72) then grbp<="011";
	end if;
	if (cc=208 and ll=73) then grbp<="011";
	end if;
	if (cc=219 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (ll=54 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=55 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=56 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=56 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<226) then grbp<="111";
	end if;
	if (ll=57 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<210) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<221) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<226) then grbp<="111";
	end if;
	if (ll=58 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=226 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=225 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=214 and ll=69) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=200 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=209 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<225) then grbp<="111";
	end if;
	if (ll=73 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

if mode="111" then

	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (cc=218 and ll=51) then grbp<="001";
	end if;
	if (cc=227 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=227 and cc<229) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (cc=203 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=226 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=54 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=54 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=226 and ll=54) then grbp<="001";
	end if;
	if (cc=229 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (ll=55 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=55 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=55) then grbp<="001";
	end if;
	if (cc=229 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=206 and ll=56) then grbp<="001";
	end if;
	if (cc=217 and ll=56) then grbp<="001";
	end if;
	if (cc=225 and ll=56) then grbp<="001";
	end if;
	if (cc=229 and ll=56) then grbp<="001";
	end if;
	if (cc=203 and ll=57) then grbp<="001";
	end if;
	if (cc=205 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=225 and ll=57) then grbp<="001";
	end if;
	if (cc=228 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=225 and ll=58) then grbp<="001";
	end if;
	if (cc=228 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=59 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=59) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=209 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<218) then grbp<="001";
	end if;
	if (ll=60 and cc>=220 and cc<223) then grbp<="001";
	end if;
	if (ll=60 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=60) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=61 and cc>=208 and cc<210) then grbp<="001";
	end if;
	if (cc=214 and ll=61) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=61 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=225 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=213 and cc<215) then grbp<="001";
	end if;
	if (ll=62 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=225 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=63) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=225 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (ll=64 and cc>=206 and cc<209) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=216 and cc<218) then grbp<="001";
	end if;
	if (ll=64 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=64) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (cc=213 and ll=65) then grbp<="001";
	end if;
	if (cc=216 and ll=65) then grbp<="001";
	end if;
	if (cc=219 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=219 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=65) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (cc=213 and ll=66) then grbp<="001";
	end if;
	if (cc=216 and ll=66) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=228 and ll=66) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (ll=67 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=67) then grbp<="001";
	end if;
	if (cc=213 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=224 and ll=67) then grbp<="001";
	end if;
	if (cc=228 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=211 and ll=68) then grbp<="001";
	end if;
	if (cc=213 and ll=68) then grbp<="001";
	end if;
	if (cc=216 and ll=68) then grbp<="001";
	end if;
	if (cc=218 and ll=68) then grbp<="001";
	end if;
	if (cc=222 and ll=68) then grbp<="001";
	end if;
	if (cc=224 and ll=68) then grbp<="001";
	end if;
	if (cc=227 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=213 and ll=69) then grbp<="001";
	end if;
	if (cc=216 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (ll=69 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=227 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=213 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (ll=70 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (ll=70 and cc>=218 and cc<220) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=227 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<211) then grbp<="001";
	end if;
	if (ll=71 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (ll=71 and cc>=224 and cc<228) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<217) then grbp<="001";
	end if;
	if (ll=72 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (ll=72 and cc>=224 and cc<227) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (ll=73 and cc>=219 and cc<221) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=206 and ll=51) then grbp<="011";
	end if;
	if (cc=228 and ll=54) then grbp<="011";
	end if;
	if (cc=217 and ll=55) then grbp<="011";
	end if;
	if (cc=226 and ll=55) then grbp<="011";
	end if;
	if (cc=204 and ll=56) then grbp<="011";
	end if;
	if (cc=207 and ll=56) then grbp<="011";
	end if;
	if (cc=202 and ll=57) then grbp<="011";
	end if;
	if (cc=211 and ll=59) then grbp<="011";
	end if;
	if (cc=220 and ll=59) then grbp<="011";
	end if;
	if (cc=208 and ll=60) then grbp<="011";
	end if;
	if (cc=210 and ll=61) then grbp<="011";
	end if;
	if (cc=204 and ll=62) then grbp<="011";
	end if;
	if (ll=62 and cc>=204 and cc<206) then grbp<="011";
	end if;
	if (cc=224 and ll=63) then grbp<="011";
	end if;
	if (cc=205 and ll=64) then grbp<="011";
	end if;
	if (cc=225 and ll=64) then grbp<="011";
	end if;
	if (cc=227 and ll=64) then grbp<="011";
	end if;
	if (cc=206 and ll=65) then grbp<="011";
	end if;
	if (cc=218 and ll=65) then grbp<="011";
	end if;
	if (cc=202 and ll=66) then grbp<="011";
	end if;
	if (cc=210 and ll=68) then grbp<="011";
	end if;
	if (cc=212 and ll=68) then grbp<="011";
	end if;
	if (cc=228 and ll=68) then grbp<="011";
	end if;
	if (cc=211 and ll=69) then grbp<="011";
	end if;
	if (ll=69 and cc>=211 and cc<213) then grbp<="011";
	end if;
	if (cc=222 and ll=70) then grbp<="011";
	end if;
	if (cc=226 and ll=70) then grbp<="011";
	end if;
	if (cc=201 and ll=73) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=203 and cc<206) then grbp<="011";
	end if;
	if (cc=213 and ll=73) then grbp<="011";
	end if;
	if (ll=73 and cc>=213 and cc<216) then grbp<="011";
	end if;
	if (cc=226 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;
	if (cc=228 and ll=78) then grbp<="011";
	end if;
	if (cc=200 and ll=79) then grbp<="011";
	end if;
	if (ll=79 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=51 and cc>=219 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=52 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=53) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=53 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=54) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<218) then grbp<="111";
	end if;
	if (ll=54 and cc>=219 and cc<226) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=55 and cc>=227 and cc<229) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=56 and cc>=226 and cc<229) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=57 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<215) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=58 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=59 and cc>=226 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (ll=60 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=61) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=212 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=61) then grbp<="111";
	end if;
	if (cc=221 and ll=61) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=61 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=209 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=215 and ll=62) then grbp<="111";
	end if;
	if (cc=218 and ll=62) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=63) then grbp<="111";
	end if;
	if (cc=209 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=220 and cc<222) then grbp<="111";
	end if;
	if (cc=229 and ll=63) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=64 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (cc=226 and ll=64) then grbp<="111";
	end if;
	if (cc=229 and ll=64) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (cc=225 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=66) then grbp<="111";
	end if;
	if (cc=225 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<224) then grbp<="111";
	end if;
	if (ll=67 and cc>=225 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=68 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<222) then grbp<="111";
	end if;
	if (cc=225 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=217 and ll=69) then grbp<="111";
	end if;
	if (cc=219 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (cc=225 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<227) then grbp<="111";
	end if;
	if (ll=69 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=70 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=217 and ll=70) then grbp<="111";
	end if;
	if (cc=220 and ll=70) then grbp<="111";
	end if;
	if (cc=223 and ll=70) then grbp<="111";
	end if;
	if (cc=225 and ll=70) then grbp<="111";
	end if;
	if (cc=228 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=211 and cc<213) then grbp<="111";
	end if;
	if (cc=222 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=204 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=72 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=72 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=206 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=206 and cc<208) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<219) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=73 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=228 and cc<230) then grbp<="111";
	end if;

end if;
if mode="110" then
	if (cc=203 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=51 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=51) then grbp<="001";
	end if;
	if (ll=51 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (ll=52 and cc>=203 and cc<205) then grbp<="001";
	end if;
	if (ll=52 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=52) then grbp<="001";
	end if;
	if (ll=52 and cc>=228 and cc<230) then grbp<="001";
	end if;
	if (cc=206 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=206 and cc<208) then grbp<="001";
	end if;
	if (cc=225 and ll=53) then grbp<="001";
	end if;
	if (ll=53 and cc>=225 and cc<228) then grbp<="001";
	end if;
	if (cc=228 and ll=53) then grbp<="001";
	end if;
	if (cc=203 and ll=54) then grbp<="001";
	end if;
	if (cc=206 and ll=54) then grbp<="001";
	end if;
	if (cc=217 and ll=54) then grbp<="001";
	end if;
	if (cc=228 and ll=54) then grbp<="001";
	end if;
	if (cc=203 and ll=55) then grbp<="001";
	end if;
	if (cc=206 and ll=55) then grbp<="001";
	end if;
	if (cc=217 and ll=55) then grbp<="001";
	end if;
	if (cc=228 and ll=55) then grbp<="001";
	end if;
	if (cc=203 and ll=56) then grbp<="001";
	end if;
	if (cc=205 and ll=56) then grbp<="001";
	end if;
	if (ll=56 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=228 and ll=56) then grbp<="001";
	end if;
	if (cc=202 and ll=57) then grbp<="001";
	end if;
	if (ll=57 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=57 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=227 and ll=57) then grbp<="001";
	end if;
	if (cc=202 and ll=58) then grbp<="001";
	end if;
	if (ll=58 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=58 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=217 and ll=58) then grbp<="001";
	end if;
	if (cc=227 and ll=58) then grbp<="001";
	end if;
	if (cc=202 and ll=59) then grbp<="001";
	end if;
	if (ll=59 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=59 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=59 and cc>=209 and cc<211) then grbp<="001";
	end if;
	if (ll=59 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=59 and cc>=220 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=60) then grbp<="001";
	end if;
	if (ll=60 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=60 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (ll=60 and cc>=208 and cc<212) then grbp<="001";
	end if;
	if (ll=60 and cc>=214 and cc<217) then grbp<="001";
	end if;
	if (ll=60 and cc>=219 and cc<222) then grbp<="001";
	end if;
	if (cc=202 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=202 and cc<204) then grbp<="001";
	end if;
	if (ll=61 and cc>=205 and cc<207) then grbp<="001";
	end if;
	if (cc=210 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=210 and cc<212) then grbp<="001";
	end if;
	if (cc=216 and ll=61) then grbp<="001";
	end if;
	if (cc=219 and ll=61) then grbp<="001";
	end if;
	if (cc=221 and ll=61) then grbp<="001";
	end if;
	if (ll=61 and cc>=221 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=62) then grbp<="001";
	end if;
	if (ll=62 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=208 and ll=62) then grbp<="001";
	end if;
	if (cc=211 and ll=62) then grbp<="001";
	end if;
	if (cc=213 and ll=62) then grbp<="001";
	end if;
	if (cc=216 and ll=62) then grbp<="001";
	end if;
	if (cc=219 and ll=62) then grbp<="001";
	end if;
	if (cc=222 and ll=62) then grbp<="001";
	end if;
	if (cc=226 and ll=62) then grbp<="001";
	end if;
	if (cc=202 and ll=63) then grbp<="001";
	end if;
	if (ll=63 and cc>=202 and cc<205) then grbp<="001";
	end if;
	if (cc=211 and ll=63) then grbp<="001";
	end if;
	if (cc=213 and ll=63) then grbp<="001";
	end if;
	if (cc=216 and ll=63) then grbp<="001";
	end if;
	if (cc=218 and ll=63) then grbp<="001";
	end if;
	if (cc=222 and ll=63) then grbp<="001";
	end if;
	if (cc=226 and ll=63) then grbp<="001";
	end if;
	if (cc=202 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=64) then grbp<="001";
	end if;
	if (cc=213 and ll=64) then grbp<="001";
	end if;
	if (cc=216 and ll=64) then grbp<="001";
	end if;
	if (cc=218 and ll=64) then grbp<="001";
	end if;
	if (ll=64 and cc>=218 and cc<223) then grbp<="001";
	end if;
	if (cc=202 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=202 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=65) then grbp<="001";
	end if;
	if (ll=65 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=66) then grbp<="001";
	end if;
	if (cc=203 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=203 and cc<206) then grbp<="001";
	end if;
	if (cc=211 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=211 and cc<213) then grbp<="001";
	end if;
	if (cc=218 and ll=66) then grbp<="001";
	end if;
	if (ll=66 and cc>=218 and cc<222) then grbp<="001";
	end if;
	if (cc=201 and ll=67) then grbp<="001";
	end if;
	if (cc=203 and ll=67) then grbp<="001";
	end if;
	if (cc=205 and ll=67) then grbp<="001";
	end if;
	if (cc=207 and ll=67) then grbp<="001";
	end if;
	if (cc=210 and ll=67) then grbp<="001";
	end if;
	if (cc=212 and ll=67) then grbp<="001";
	end if;
	if (cc=216 and ll=67) then grbp<="001";
	end if;
	if (cc=218 and ll=67) then grbp<="001";
	end if;
	if (cc=225 and ll=67) then grbp<="001";
	end if;
	if (cc=201 and ll=68) then grbp<="001";
	end if;
	if (cc=203 and ll=68) then grbp<="001";
	end if;
	if (cc=205 and ll=68) then grbp<="001";
	end if;
	if (cc=207 and ll=68) then grbp<="001";
	end if;
	if (cc=210 and ll=68) then grbp<="001";
	end if;
	if (cc=212 and ll=68) then grbp<="001";
	end if;
	if (cc=215 and ll=68) then grbp<="001";
	end if;
	if (ll=68 and cc>=215 and cc<217) then grbp<="001";
	end if;
	if (cc=221 and ll=68) then grbp<="001";
	end if;
	if (cc=225 and ll=68) then grbp<="001";
	end if;
	if (cc=201 and ll=69) then grbp<="001";
	end if;
	if (cc=203 and ll=69) then grbp<="001";
	end if;
	if (cc=205 and ll=69) then grbp<="001";
	end if;
	if (cc=207 and ll=69) then grbp<="001";
	end if;
	if (cc=210 and ll=69) then grbp<="001";
	end if;
	if (cc=212 and ll=69) then grbp<="001";
	end if;
	if (cc=215 and ll=69) then grbp<="001";
	end if;
	if (cc=218 and ll=69) then grbp<="001";
	end if;
	if (cc=221 and ll=69) then grbp<="001";
	end if;
	if (cc=224 and ll=69) then grbp<="001";
	end if;
	if (cc=201 and ll=70) then grbp<="001";
	end if;
	if (cc=203 and ll=70) then grbp<="001";
	end if;
	if (cc=205 and ll=70) then grbp<="001";
	end if;
	if (cc=207 and ll=70) then grbp<="001";
	end if;
	if (cc=210 and ll=70) then grbp<="001";
	end if;
	if (cc=212 and ll=70) then grbp<="001";
	end if;
	if (cc=215 and ll=70) then grbp<="001";
	end if;
	if (cc=218 and ll=70) then grbp<="001";
	end if;
	if (cc=221 and ll=70) then grbp<="001";
	end if;
	if (cc=224 and ll=70) then grbp<="001";
	end if;
	if (cc=201 and ll=71) then grbp<="001";
	end if;
	if (cc=203 and ll=71) then grbp<="001";
	end if;
	if (cc=205 and ll=71) then grbp<="001";
	end if;
	if (cc=207 and ll=71) then grbp<="001";
	end if;
	if (ll=71 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=71 and cc>=212 and cc<216) then grbp<="001";
	end if;
	if (ll=71 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=72) then grbp<="001";
	end if;
	if (cc=203 and ll=72) then grbp<="001";
	end if;
	if (cc=205 and ll=72) then grbp<="001";
	end if;
	if (cc=207 and ll=72) then grbp<="001";
	end if;
	if (ll=72 and cc>=207 and cc<210) then grbp<="001";
	end if;
	if (ll=72 and cc>=213 and cc<216) then grbp<="001";
	end if;
	if (ll=72 and cc>=218 and cc<221) then grbp<="001";
	end if;
	if (cc=201 and ll=73) then grbp<="001";
	end if;
	if (cc=204 and ll=73) then grbp<="001";
	end if;
	if (cc=208 and ll=73) then grbp<="001";
	end if;
	if (cc=213 and ll=73) then grbp<="001";
	end if;
	if (cc=215 and ll=73) then grbp<="001";
	end if;
	if (cc=219 and ll=73) then grbp<="001";
	end if;
	if (cc=224 and ll=73) then grbp<="001";
	end if;
	if (cc=200 and ll=78) then grbp<="001";
	end if;
	if (ll=78 and cc>=200 and cc<228) then grbp<="001";
	end if;

	if (cc=229 and ll=53) then grbp<="011";
	end if;
	if (cc=207 and ll=54) then grbp<="011";
	end if;
	if (cc=202 and ll=56) then grbp<="011";
	end if;
	if (cc=227 and ll=56) then grbp<="011";
	end if;
	if (cc=209 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=209 and cc<211) then grbp<="011";
	end if;
	if (cc=220 and ll=58) then grbp<="011";
	end if;
	if (ll=58 and cc>=220 and cc<222) then grbp<="011";
	end if;
	if (cc=213 and ll=60) then grbp<="011";
	end if;
	if (cc=222 and ll=60) then grbp<="011";
	end if;
	if (cc=227 and ll=60) then grbp<="011";
	end if;
	if (cc=204 and ll=61) then grbp<="011";
	end if;
	if (cc=209 and ll=61) then grbp<="011";
	end if;
	if (cc=214 and ll=61) then grbp<="011";
	end if;
	if (cc=205 and ll=62) then grbp<="011";
	end if;
	if (cc=207 and ll=62) then grbp<="011";
	end if;
	if (cc=218 and ll=62) then grbp<="011";
	end if;
	if (cc=221 and ll=62) then grbp<="011";
	end if;
	if (cc=205 and ll=63) then grbp<="011";
	end if;
	if (ll=63 and cc>=205 and cc<207) then grbp<="011";
	end if;
	if (cc=221 and ll=63) then grbp<="011";
	end if;
	if (cc=226 and ll=64) then grbp<="011";
	end if;
	if (cc=201 and ll=65) then grbp<="011";
	end if;
	if (cc=213 and ll=65) then grbp<="011";
	end if;
	if (cc=222 and ll=65) then grbp<="011";
	end if;
	if (cc=210 and ll=66) then grbp<="011";
	end if;
	if (cc=204 and ll=67) then grbp<="011";
	end if;
	if (cc=211 and ll=67) then grbp<="011";
	end if;
	if (cc=224 and ll=68) then grbp<="011";
	end if;
	if (cc=209 and ll=70) then grbp<="011";
	end if;
	if (cc=213 and ll=70) then grbp<="011";
	end if;
	if (cc=220 and ll=70) then grbp<="011";
	end if;
	if (cc=210 and ll=71) then grbp<="011";
	end if;
	if (cc=221 and ll=71) then grbp<="011";
	end if;
	if (cc=204 and ll=72) then grbp<="011";
	end if;
	if (cc=212 and ll=72) then grbp<="011";
	end if;
	if (cc=203 and ll=73) then grbp<="011";
	end if;
	if (cc=207 and ll=73) then grbp<="011";
	end if;
	if (cc=209 and ll=73) then grbp<="011";
	end if;
	if (cc=214 and ll=73) then grbp<="011";
	end if;
	if (cc=218 and ll=73) then grbp<="011";
	end if;
	if (cc=220 and ll=73) then grbp<="011";
	end if;
	if (cc=223 and ll=73) then grbp<="011";
	end if;
	if (cc=200 and ll=77) then grbp<="011";
	end if;
	if (ll=77 and cc>=200 and cc<228) then grbp<="011";
	end if;


	if (cc=200 and ll=50) then grbp<="111";
	end if;
	if (ll=50 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=51) then grbp<="111";
	end if;
	if (ll=51 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=51 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=52 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (cc=208 and ll=52) then grbp<="111";
	end if;
	if (ll=52 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=52 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=53 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=53 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=53 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=53 and cc>=218 and cc<225) then grbp<="111";
	end if;
	if (ll=54 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=54 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=54 and cc>=208 and cc<217) then grbp<="111";
	end if;
	if (ll=54 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=55) then grbp<="111";
	end if;
	if (ll=55 and cc>=200 and cc<203) then grbp<="111";
	end if;
	if (ll=55 and cc>=204 and cc<206) then grbp<="111";
	end if;
	if (ll=55 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=55 and cc>=218 and cc<228) then grbp<="111";
	end if;
	if (cc=200 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=56) then grbp<="111";
	end if;
	if (ll=56 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=56 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (cc=200 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=57) then grbp<="111";
	end if;
	if (ll=57 and cc>=207 and cc<217) then grbp<="111";
	end if;
	if (ll=57 and cc>=218 and cc<227) then grbp<="111";
	end if;
	if (ll=57 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=58 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (cc=218 and ll=58) then grbp<="111";
	end if;
	if (ll=58 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=58 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=58 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=59) then grbp<="111";
	end if;
	if (ll=59 and cc>=207 and cc<209) then grbp<="111";
	end if;
	if (ll=59 and cc>=211 and cc<214) then grbp<="111";
	end if;
	if (ll=59 and cc>=218 and cc<220) then grbp<="111";
	end if;
	if (ll=59 and cc>=222 and cc<227) then grbp<="111";
	end if;
	if (ll=59 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=207 and ll=60) then grbp<="111";
	end if;
	if (cc=212 and ll=60) then grbp<="111";
	end if;
	if (cc=217 and ll=60) then grbp<="111";
	end if;
	if (ll=60 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (ll=60 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=60 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=212 and ll=61) then grbp<="111";
	end if;
	if (cc=215 and ll=61) then grbp<="111";
	end if;
	if (cc=217 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=217 and cc<219) then grbp<="111";
	end if;
	if (cc=223 and ll=61) then grbp<="111";
	end if;
	if (ll=61 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=61 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=62 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=220 and ll=62) then grbp<="111";
	end if;
	if (cc=223 and ll=62) then grbp<="111";
	end if;
	if (ll=62 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=62 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (ll=63 and cc>=209 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=63) then grbp<="111";
	end if;
	if (ll=63 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=63 and cc>=223 and cc<226) then grbp<="111";
	end if;
	if (ll=63 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=200 and cc<202) then grbp<="111";
	end if;
	if (cc=208 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (cc=214 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=64) then grbp<="111";
	end if;
	if (ll=64 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=64 and cc>=227 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=65) then grbp<="111";
	end if;
	if (cc=206 and ll=65) then grbp<="111";
	end if;
	if (cc=208 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=208 and cc<211) then grbp<="111";
	end if;
	if (ll=65 and cc>=214 and cc<216) then grbp<="111";
	end if;
	if (cc=223 and ll=65) then grbp<="111";
	end if;
	if (ll=65 and cc>=223 and cc<225) then grbp<="111";
	end if;
	if (ll=65 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=66) then grbp<="111";
	end if;
	if (cc=202 and ll=66) then grbp<="111";
	end if;
	if (cc=206 and ll=66) then grbp<="111";
	end if;
	if (cc=208 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=66 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=222 and ll=66) then grbp<="111";
	end if;
	if (ll=66 and cc>=222 and cc<225) then grbp<="111";
	end if;
	if (ll=66 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=67) then grbp<="111";
	end if;
	if (cc=202 and ll=67) then grbp<="111";
	end if;
	if (cc=206 and ll=67) then grbp<="111";
	end if;
	if (cc=208 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (ll=67 and cc>=213 and cc<216) then grbp<="111";
	end if;
	if (cc=219 and ll=67) then grbp<="111";
	end if;
	if (ll=67 and cc>=219 and cc<225) then grbp<="111";
	end if;
	if (ll=67 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=68) then grbp<="111";
	end if;
	if (cc=202 and ll=68) then grbp<="111";
	end if;
	if (cc=204 and ll=68) then grbp<="111";
	end if;
	if (cc=206 and ll=68) then grbp<="111";
	end if;
	if (cc=208 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (cc=219 and ll=68) then grbp<="111";
	end if;
	if (ll=68 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=68 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=68 and cc>=226 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=69) then grbp<="111";
	end if;
	if (cc=202 and ll=69) then grbp<="111";
	end if;
	if (cc=204 and ll=69) then grbp<="111";
	end if;
	if (cc=206 and ll=69) then grbp<="111";
	end if;
	if (cc=208 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=208 and cc<210) then grbp<="111";
	end if;
	if (cc=213 and ll=69) then grbp<="111";
	end if;
	if (ll=69 and cc>=213 and cc<215) then grbp<="111";
	end if;
	if (ll=69 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=69 and cc>=219 and cc<221) then grbp<="111";
	end if;
	if (ll=69 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=69 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=70) then grbp<="111";
	end if;
	if (cc=202 and ll=70) then grbp<="111";
	end if;
	if (cc=204 and ll=70) then grbp<="111";
	end if;
	if (cc=206 and ll=70) then grbp<="111";
	end if;
	if (cc=208 and ll=70) then grbp<="111";
	end if;
	if (cc=211 and ll=70) then grbp<="111";
	end if;
	if (cc=214 and ll=70) then grbp<="111";
	end if;
	if (cc=216 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (cc=222 and ll=70) then grbp<="111";
	end if;
	if (ll=70 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=70 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=71) then grbp<="111";
	end if;
	if (cc=202 and ll=71) then grbp<="111";
	end if;
	if (cc=204 and ll=71) then grbp<="111";
	end if;
	if (cc=206 and ll=71) then grbp<="111";
	end if;
	if (cc=211 and ll=71) then grbp<="111";
	end if;
	if (cc=216 and ll=71) then grbp<="111";
	end if;
	if (ll=71 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=71 and cc>=222 and cc<224) then grbp<="111";
	end if;
	if (ll=71 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=72) then grbp<="111";
	end if;
	if (cc=202 and ll=72) then grbp<="111";
	end if;
	if (cc=206 and ll=72) then grbp<="111";
	end if;
	if (cc=210 and ll=72) then grbp<="111";
	end if;
	if (ll=72 and cc>=210 and cc<212) then grbp<="111";
	end if;
	if (ll=72 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=72 and cc>=221 and cc<224) then grbp<="111";
	end if;
	if (ll=72 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=73) then grbp<="111";
	end if;
	if (cc=202 and ll=73) then grbp<="111";
	end if;
	if (cc=205 and ll=73) then grbp<="111";
	end if;
	if (ll=73 and cc>=205 and cc<207) then grbp<="111";
	end if;
	if (ll=73 and cc>=210 and cc<213) then grbp<="111";
	end if;
	if (ll=73 and cc>=216 and cc<218) then grbp<="111";
	end if;
	if (ll=73 and cc>=221 and cc<223) then grbp<="111";
	end if;
	if (ll=73 and cc>=225 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=74) then grbp<="111";
	end if;
	if (ll=74 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=75) then grbp<="111";
	end if;
	if (ll=75 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=76) then grbp<="111";
	end if;
	if (ll=76 and cc>=200 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=77) then grbp<="111";
	end if;
	if (ll=77 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=228 and ll=78) then grbp<="111";
	end if;
	if (ll=78 and cc>=228 and cc<230) then grbp<="111";
	end if;
	if (cc=200 and ll=79) then grbp<="111";
	end if;
	if (ll=79 and cc>=200 and cc<230) then grbp<="111";
	end if;

end if;

end process;

hs<=hs1;vs<=vs1;r<=grb(2);g<=grb(3);b<=grb(1);

end one;
